import MemTypes::*;
import ProcTypes::*;

// Python generated code which returns arc_id for each pair of source and destination of packets 

function NoCArcId lookupNoCArcId(ProcID srcProcId, ProcID destProcID);
  if (srcProcId == 0) begin
    if(destProcID == 1) return 0;
    if(destProcID == 3) return 1;
    if(destProcID == 12) return 2;
    if(destProcID == 20) return 3;
    if(destProcID == 34) return 4;
    if(destProcID == 38) return 5;
    if(destProcID == 81) return 6;
    if(destProcID == 88) return 7;
    if(destProcID == 94) return 8;
    if(destProcID == 104) return 9;
    if(destProcID == 109) return 10;
    if(destProcID == 132) return 11;
    if(destProcID == 130) return 12;
    if(destProcID == 121) return 13;
    if(destProcID == 113) return 14;
    if(destProcID == 99) return 15;
    if(destProcID == 95) return 16;
    if(destProcID == 52) return 17;
    if(destProcID == 45) return 18;
    if(destProcID == 39) return 19;
    if(destProcID == 29) return 20;
    if(destProcID == 24) return 21;
  end
  if (srcProcId == 1) begin
    if(destProcID == 2) return 22;
    if(destProcID == 4) return 23;
    if(destProcID == 13) return 24;
    if(destProcID == 21) return 25;
    if(destProcID == 35) return 26;
    if(destProcID == 39) return 27;
    if(destProcID == 82) return 28;
    if(destProcID == 89) return 29;
    if(destProcID == 95) return 30;
    if(destProcID == 105) return 31;
    if(destProcID == 110) return 32;
    if(destProcID == 0) return 33;
    if(destProcID == 131) return 34;
    if(destProcID == 122) return 35;
    if(destProcID == 114) return 36;
    if(destProcID == 100) return 37;
    if(destProcID == 96) return 38;
    if(destProcID == 53) return 39;
    if(destProcID == 46) return 40;
    if(destProcID == 40) return 41;
    if(destProcID == 30) return 42;
    if(destProcID == 25) return 43;
  end
  if (srcProcId == 2) begin
    if(destProcID == 3) return 44;
    if(destProcID == 5) return 45;
    if(destProcID == 14) return 46;
    if(destProcID == 22) return 47;
    if(destProcID == 36) return 48;
    if(destProcID == 40) return 49;
    if(destProcID == 83) return 50;
    if(destProcID == 90) return 51;
    if(destProcID == 96) return 52;
    if(destProcID == 106) return 53;
    if(destProcID == 111) return 54;
    if(destProcID == 1) return 55;
    if(destProcID == 132) return 56;
    if(destProcID == 123) return 57;
    if(destProcID == 115) return 58;
    if(destProcID == 101) return 59;
    if(destProcID == 97) return 60;
    if(destProcID == 54) return 61;
    if(destProcID == 47) return 62;
    if(destProcID == 41) return 63;
    if(destProcID == 31) return 64;
    if(destProcID == 26) return 65;
  end
  if (srcProcId == 3) begin
    if(destProcID == 4) return 66;
    if(destProcID == 6) return 67;
    if(destProcID == 15) return 68;
    if(destProcID == 23) return 69;
    if(destProcID == 37) return 70;
    if(destProcID == 41) return 71;
    if(destProcID == 84) return 72;
    if(destProcID == 91) return 73;
    if(destProcID == 97) return 74;
    if(destProcID == 107) return 75;
    if(destProcID == 112) return 76;
    if(destProcID == 2) return 77;
    if(destProcID == 0) return 78;
    if(destProcID == 124) return 79;
    if(destProcID == 116) return 80;
    if(destProcID == 102) return 81;
    if(destProcID == 98) return 82;
    if(destProcID == 55) return 83;
    if(destProcID == 48) return 84;
    if(destProcID == 42) return 85;
    if(destProcID == 32) return 86;
    if(destProcID == 27) return 87;
  end
  if (srcProcId == 4) begin
    if(destProcID == 5) return 88;
    if(destProcID == 7) return 89;
    if(destProcID == 16) return 90;
    if(destProcID == 24) return 91;
    if(destProcID == 38) return 92;
    if(destProcID == 42) return 93;
    if(destProcID == 85) return 94;
    if(destProcID == 92) return 95;
    if(destProcID == 98) return 96;
    if(destProcID == 108) return 97;
    if(destProcID == 113) return 98;
    if(destProcID == 3) return 99;
    if(destProcID == 1) return 100;
    if(destProcID == 125) return 101;
    if(destProcID == 117) return 102;
    if(destProcID == 103) return 103;
    if(destProcID == 99) return 104;
    if(destProcID == 56) return 105;
    if(destProcID == 49) return 106;
    if(destProcID == 43) return 107;
    if(destProcID == 33) return 108;
    if(destProcID == 28) return 109;
  end
  if (srcProcId == 5) begin
    if(destProcID == 6) return 110;
    if(destProcID == 8) return 111;
    if(destProcID == 17) return 112;
    if(destProcID == 25) return 113;
    if(destProcID == 39) return 114;
    if(destProcID == 43) return 115;
    if(destProcID == 86) return 116;
    if(destProcID == 93) return 117;
    if(destProcID == 99) return 118;
    if(destProcID == 109) return 119;
    if(destProcID == 114) return 120;
    if(destProcID == 4) return 121;
    if(destProcID == 2) return 122;
    if(destProcID == 126) return 123;
    if(destProcID == 118) return 124;
    if(destProcID == 104) return 125;
    if(destProcID == 100) return 126;
    if(destProcID == 57) return 127;
    if(destProcID == 50) return 128;
    if(destProcID == 44) return 129;
    if(destProcID == 34) return 130;
    if(destProcID == 29) return 131;
  end
  if (srcProcId == 6) begin
    if(destProcID == 7) return 132;
    if(destProcID == 9) return 133;
    if(destProcID == 18) return 134;
    if(destProcID == 26) return 135;
    if(destProcID == 40) return 136;
    if(destProcID == 44) return 137;
    if(destProcID == 87) return 138;
    if(destProcID == 94) return 139;
    if(destProcID == 100) return 140;
    if(destProcID == 110) return 141;
    if(destProcID == 115) return 142;
    if(destProcID == 5) return 143;
    if(destProcID == 3) return 144;
    if(destProcID == 127) return 145;
    if(destProcID == 119) return 146;
    if(destProcID == 105) return 147;
    if(destProcID == 101) return 148;
    if(destProcID == 58) return 149;
    if(destProcID == 51) return 150;
    if(destProcID == 45) return 151;
    if(destProcID == 35) return 152;
    if(destProcID == 30) return 153;
  end
  if (srcProcId == 7) begin
    if(destProcID == 8) return 154;
    if(destProcID == 10) return 155;
    if(destProcID == 19) return 156;
    if(destProcID == 27) return 157;
    if(destProcID == 41) return 158;
    if(destProcID == 45) return 159;
    if(destProcID == 88) return 160;
    if(destProcID == 95) return 161;
    if(destProcID == 101) return 162;
    if(destProcID == 111) return 163;
    if(destProcID == 116) return 164;
    if(destProcID == 6) return 165;
    if(destProcID == 4) return 166;
    if(destProcID == 128) return 167;
    if(destProcID == 120) return 168;
    if(destProcID == 106) return 169;
    if(destProcID == 102) return 170;
    if(destProcID == 59) return 171;
    if(destProcID == 52) return 172;
    if(destProcID == 46) return 173;
    if(destProcID == 36) return 174;
    if(destProcID == 31) return 175;
  end
  if (srcProcId == 8) begin
    if(destProcID == 9) return 176;
    if(destProcID == 11) return 177;
    if(destProcID == 20) return 178;
    if(destProcID == 28) return 179;
    if(destProcID == 42) return 180;
    if(destProcID == 46) return 181;
    if(destProcID == 89) return 182;
    if(destProcID == 96) return 183;
    if(destProcID == 102) return 184;
    if(destProcID == 112) return 185;
    if(destProcID == 117) return 186;
    if(destProcID == 7) return 187;
    if(destProcID == 5) return 188;
    if(destProcID == 129) return 189;
    if(destProcID == 121) return 190;
    if(destProcID == 107) return 191;
    if(destProcID == 103) return 192;
    if(destProcID == 60) return 193;
    if(destProcID == 53) return 194;
    if(destProcID == 47) return 195;
    if(destProcID == 37) return 196;
    if(destProcID == 32) return 197;
  end
  if (srcProcId == 9) begin
    if(destProcID == 10) return 198;
    if(destProcID == 12) return 199;
    if(destProcID == 21) return 200;
    if(destProcID == 29) return 201;
    if(destProcID == 43) return 202;
    if(destProcID == 47) return 203;
    if(destProcID == 90) return 204;
    if(destProcID == 97) return 205;
    if(destProcID == 103) return 206;
    if(destProcID == 113) return 207;
    if(destProcID == 118) return 208;
    if(destProcID == 8) return 209;
    if(destProcID == 6) return 210;
    if(destProcID == 130) return 211;
    if(destProcID == 122) return 212;
    if(destProcID == 108) return 213;
    if(destProcID == 104) return 214;
    if(destProcID == 61) return 215;
    if(destProcID == 54) return 216;
    if(destProcID == 48) return 217;
    if(destProcID == 38) return 218;
    if(destProcID == 33) return 219;
  end
  if (srcProcId == 10) begin
    if(destProcID == 11) return 220;
    if(destProcID == 13) return 221;
    if(destProcID == 22) return 222;
    if(destProcID == 30) return 223;
    if(destProcID == 44) return 224;
    if(destProcID == 48) return 225;
    if(destProcID == 91) return 226;
    if(destProcID == 98) return 227;
    if(destProcID == 104) return 228;
    if(destProcID == 114) return 229;
    if(destProcID == 119) return 230;
    if(destProcID == 9) return 231;
    if(destProcID == 7) return 232;
    if(destProcID == 131) return 233;
    if(destProcID == 123) return 234;
    if(destProcID == 109) return 235;
    if(destProcID == 105) return 236;
    if(destProcID == 62) return 237;
    if(destProcID == 55) return 238;
    if(destProcID == 49) return 239;
    if(destProcID == 39) return 240;
    if(destProcID == 34) return 241;
  end
  if (srcProcId == 11) begin
    if(destProcID == 12) return 242;
    if(destProcID == 14) return 243;
    if(destProcID == 23) return 244;
    if(destProcID == 31) return 245;
    if(destProcID == 45) return 246;
    if(destProcID == 49) return 247;
    if(destProcID == 92) return 248;
    if(destProcID == 99) return 249;
    if(destProcID == 105) return 250;
    if(destProcID == 115) return 251;
    if(destProcID == 120) return 252;
    if(destProcID == 10) return 253;
    if(destProcID == 8) return 254;
    if(destProcID == 132) return 255;
    if(destProcID == 124) return 256;
    if(destProcID == 110) return 257;
    if(destProcID == 106) return 258;
    if(destProcID == 63) return 259;
    if(destProcID == 56) return 260;
    if(destProcID == 50) return 261;
    if(destProcID == 40) return 262;
    if(destProcID == 35) return 263;
  end
  if (srcProcId == 12) begin
    if(destProcID == 13) return 264;
    if(destProcID == 15) return 265;
    if(destProcID == 24) return 266;
    if(destProcID == 32) return 267;
    if(destProcID == 46) return 268;
    if(destProcID == 50) return 269;
    if(destProcID == 93) return 270;
    if(destProcID == 100) return 271;
    if(destProcID == 106) return 272;
    if(destProcID == 116) return 273;
    if(destProcID == 121) return 274;
    if(destProcID == 11) return 275;
    if(destProcID == 9) return 276;
    if(destProcID == 0) return 277;
    if(destProcID == 125) return 278;
    if(destProcID == 111) return 279;
    if(destProcID == 107) return 280;
    if(destProcID == 64) return 281;
    if(destProcID == 57) return 282;
    if(destProcID == 51) return 283;
    if(destProcID == 41) return 284;
    if(destProcID == 36) return 285;
  end
  if (srcProcId == 13) begin
    if(destProcID == 14) return 286;
    if(destProcID == 16) return 287;
    if(destProcID == 25) return 288;
    if(destProcID == 33) return 289;
    if(destProcID == 47) return 290;
    if(destProcID == 51) return 291;
    if(destProcID == 94) return 292;
    if(destProcID == 101) return 293;
    if(destProcID == 107) return 294;
    if(destProcID == 117) return 295;
    if(destProcID == 122) return 296;
    if(destProcID == 12) return 297;
    if(destProcID == 10) return 298;
    if(destProcID == 1) return 299;
    if(destProcID == 126) return 300;
    if(destProcID == 112) return 301;
    if(destProcID == 108) return 302;
    if(destProcID == 65) return 303;
    if(destProcID == 58) return 304;
    if(destProcID == 52) return 305;
    if(destProcID == 42) return 306;
    if(destProcID == 37) return 307;
  end
  if (srcProcId == 14) begin
    if(destProcID == 15) return 308;
    if(destProcID == 17) return 309;
    if(destProcID == 26) return 310;
    if(destProcID == 34) return 311;
    if(destProcID == 48) return 312;
    if(destProcID == 52) return 313;
    if(destProcID == 95) return 314;
    if(destProcID == 102) return 315;
    if(destProcID == 108) return 316;
    if(destProcID == 118) return 317;
    if(destProcID == 123) return 318;
    if(destProcID == 13) return 319;
    if(destProcID == 11) return 320;
    if(destProcID == 2) return 321;
    if(destProcID == 127) return 322;
    if(destProcID == 113) return 323;
    if(destProcID == 109) return 324;
    if(destProcID == 66) return 325;
    if(destProcID == 59) return 326;
    if(destProcID == 53) return 327;
    if(destProcID == 43) return 328;
    if(destProcID == 38) return 329;
  end
  if (srcProcId == 15) begin
    if(destProcID == 16) return 330;
    if(destProcID == 18) return 331;
    if(destProcID == 27) return 332;
    if(destProcID == 35) return 333;
    if(destProcID == 49) return 334;
    if(destProcID == 53) return 335;
    if(destProcID == 96) return 336;
    if(destProcID == 103) return 337;
    if(destProcID == 109) return 338;
    if(destProcID == 119) return 339;
    if(destProcID == 124) return 340;
    if(destProcID == 14) return 341;
    if(destProcID == 12) return 342;
    if(destProcID == 3) return 343;
    if(destProcID == 128) return 344;
    if(destProcID == 114) return 345;
    if(destProcID == 110) return 346;
    if(destProcID == 67) return 347;
    if(destProcID == 60) return 348;
    if(destProcID == 54) return 349;
    if(destProcID == 44) return 350;
    if(destProcID == 39) return 351;
  end
  if (srcProcId == 16) begin
    if(destProcID == 17) return 352;
    if(destProcID == 19) return 353;
    if(destProcID == 28) return 354;
    if(destProcID == 36) return 355;
    if(destProcID == 50) return 356;
    if(destProcID == 54) return 357;
    if(destProcID == 97) return 358;
    if(destProcID == 104) return 359;
    if(destProcID == 110) return 360;
    if(destProcID == 120) return 361;
    if(destProcID == 125) return 362;
    if(destProcID == 15) return 363;
    if(destProcID == 13) return 364;
    if(destProcID == 4) return 365;
    if(destProcID == 129) return 366;
    if(destProcID == 115) return 367;
    if(destProcID == 111) return 368;
    if(destProcID == 68) return 369;
    if(destProcID == 61) return 370;
    if(destProcID == 55) return 371;
    if(destProcID == 45) return 372;
    if(destProcID == 40) return 373;
  end
  if (srcProcId == 17) begin
    if(destProcID == 18) return 374;
    if(destProcID == 20) return 375;
    if(destProcID == 29) return 376;
    if(destProcID == 37) return 377;
    if(destProcID == 51) return 378;
    if(destProcID == 55) return 379;
    if(destProcID == 98) return 380;
    if(destProcID == 105) return 381;
    if(destProcID == 111) return 382;
    if(destProcID == 121) return 383;
    if(destProcID == 126) return 384;
    if(destProcID == 16) return 385;
    if(destProcID == 14) return 386;
    if(destProcID == 5) return 387;
    if(destProcID == 130) return 388;
    if(destProcID == 116) return 389;
    if(destProcID == 112) return 390;
    if(destProcID == 69) return 391;
    if(destProcID == 62) return 392;
    if(destProcID == 56) return 393;
    if(destProcID == 46) return 394;
    if(destProcID == 41) return 395;
  end
  if (srcProcId == 18) begin
    if(destProcID == 19) return 396;
    if(destProcID == 21) return 397;
    if(destProcID == 30) return 398;
    if(destProcID == 38) return 399;
    if(destProcID == 52) return 400;
    if(destProcID == 56) return 401;
    if(destProcID == 99) return 402;
    if(destProcID == 106) return 403;
    if(destProcID == 112) return 404;
    if(destProcID == 122) return 405;
    if(destProcID == 127) return 406;
    if(destProcID == 17) return 407;
    if(destProcID == 15) return 408;
    if(destProcID == 6) return 409;
    if(destProcID == 131) return 410;
    if(destProcID == 117) return 411;
    if(destProcID == 113) return 412;
    if(destProcID == 70) return 413;
    if(destProcID == 63) return 414;
    if(destProcID == 57) return 415;
    if(destProcID == 47) return 416;
    if(destProcID == 42) return 417;
  end
  if (srcProcId == 19) begin
    if(destProcID == 20) return 418;
    if(destProcID == 22) return 419;
    if(destProcID == 31) return 420;
    if(destProcID == 39) return 421;
    if(destProcID == 53) return 422;
    if(destProcID == 57) return 423;
    if(destProcID == 100) return 424;
    if(destProcID == 107) return 425;
    if(destProcID == 113) return 426;
    if(destProcID == 123) return 427;
    if(destProcID == 128) return 428;
    if(destProcID == 18) return 429;
    if(destProcID == 16) return 430;
    if(destProcID == 7) return 431;
    if(destProcID == 132) return 432;
    if(destProcID == 118) return 433;
    if(destProcID == 114) return 434;
    if(destProcID == 71) return 435;
    if(destProcID == 64) return 436;
    if(destProcID == 58) return 437;
    if(destProcID == 48) return 438;
    if(destProcID == 43) return 439;
  end
  if (srcProcId == 20) begin
    if(destProcID == 21) return 440;
    if(destProcID == 23) return 441;
    if(destProcID == 32) return 442;
    if(destProcID == 40) return 443;
    if(destProcID == 54) return 444;
    if(destProcID == 58) return 445;
    if(destProcID == 101) return 446;
    if(destProcID == 108) return 447;
    if(destProcID == 114) return 448;
    if(destProcID == 124) return 449;
    if(destProcID == 129) return 450;
    if(destProcID == 19) return 451;
    if(destProcID == 17) return 452;
    if(destProcID == 8) return 453;
    if(destProcID == 0) return 454;
    if(destProcID == 119) return 455;
    if(destProcID == 115) return 456;
    if(destProcID == 72) return 457;
    if(destProcID == 65) return 458;
    if(destProcID == 59) return 459;
    if(destProcID == 49) return 460;
    if(destProcID == 44) return 461;
  end
  if (srcProcId == 21) begin
    if(destProcID == 22) return 462;
    if(destProcID == 24) return 463;
    if(destProcID == 33) return 464;
    if(destProcID == 41) return 465;
    if(destProcID == 55) return 466;
    if(destProcID == 59) return 467;
    if(destProcID == 102) return 468;
    if(destProcID == 109) return 469;
    if(destProcID == 115) return 470;
    if(destProcID == 125) return 471;
    if(destProcID == 130) return 472;
    if(destProcID == 20) return 473;
    if(destProcID == 18) return 474;
    if(destProcID == 9) return 475;
    if(destProcID == 1) return 476;
    if(destProcID == 120) return 477;
    if(destProcID == 116) return 478;
    if(destProcID == 73) return 479;
    if(destProcID == 66) return 480;
    if(destProcID == 60) return 481;
    if(destProcID == 50) return 482;
    if(destProcID == 45) return 483;
  end
  if (srcProcId == 22) begin
    if(destProcID == 23) return 484;
    if(destProcID == 25) return 485;
    if(destProcID == 34) return 486;
    if(destProcID == 42) return 487;
    if(destProcID == 56) return 488;
    if(destProcID == 60) return 489;
    if(destProcID == 103) return 490;
    if(destProcID == 110) return 491;
    if(destProcID == 116) return 492;
    if(destProcID == 126) return 493;
    if(destProcID == 131) return 494;
    if(destProcID == 21) return 495;
    if(destProcID == 19) return 496;
    if(destProcID == 10) return 497;
    if(destProcID == 2) return 498;
    if(destProcID == 121) return 499;
    if(destProcID == 117) return 500;
    if(destProcID == 74) return 501;
    if(destProcID == 67) return 502;
    if(destProcID == 61) return 503;
    if(destProcID == 51) return 504;
    if(destProcID == 46) return 505;
  end
  if (srcProcId == 23) begin
    if(destProcID == 24) return 506;
    if(destProcID == 26) return 507;
    if(destProcID == 35) return 508;
    if(destProcID == 43) return 509;
    if(destProcID == 57) return 510;
    if(destProcID == 61) return 511;
    if(destProcID == 104) return 512;
    if(destProcID == 111) return 513;
    if(destProcID == 117) return 514;
    if(destProcID == 127) return 515;
    if(destProcID == 132) return 516;
    if(destProcID == 22) return 517;
    if(destProcID == 20) return 518;
    if(destProcID == 11) return 519;
    if(destProcID == 3) return 520;
    if(destProcID == 122) return 521;
    if(destProcID == 118) return 522;
    if(destProcID == 75) return 523;
    if(destProcID == 68) return 524;
    if(destProcID == 62) return 525;
    if(destProcID == 52) return 526;
    if(destProcID == 47) return 527;
  end
  if (srcProcId == 24) begin
    if(destProcID == 25) return 528;
    if(destProcID == 27) return 529;
    if(destProcID == 36) return 530;
    if(destProcID == 44) return 531;
    if(destProcID == 58) return 532;
    if(destProcID == 62) return 533;
    if(destProcID == 105) return 534;
    if(destProcID == 112) return 535;
    if(destProcID == 118) return 536;
    if(destProcID == 128) return 537;
    if(destProcID == 0) return 538;
    if(destProcID == 23) return 539;
    if(destProcID == 21) return 540;
    if(destProcID == 12) return 541;
    if(destProcID == 4) return 542;
    if(destProcID == 123) return 543;
    if(destProcID == 119) return 544;
    if(destProcID == 76) return 545;
    if(destProcID == 69) return 546;
    if(destProcID == 63) return 547;
    if(destProcID == 53) return 548;
    if(destProcID == 48) return 549;
  end
  if (srcProcId == 25) begin
    if(destProcID == 26) return 550;
    if(destProcID == 28) return 551;
    if(destProcID == 37) return 552;
    if(destProcID == 45) return 553;
    if(destProcID == 59) return 554;
    if(destProcID == 63) return 555;
    if(destProcID == 106) return 556;
    if(destProcID == 113) return 557;
    if(destProcID == 119) return 558;
    if(destProcID == 129) return 559;
    if(destProcID == 1) return 560;
    if(destProcID == 24) return 561;
    if(destProcID == 22) return 562;
    if(destProcID == 13) return 563;
    if(destProcID == 5) return 564;
    if(destProcID == 124) return 565;
    if(destProcID == 120) return 566;
    if(destProcID == 77) return 567;
    if(destProcID == 70) return 568;
    if(destProcID == 64) return 569;
    if(destProcID == 54) return 570;
    if(destProcID == 49) return 571;
  end
  if (srcProcId == 26) begin
    if(destProcID == 27) return 572;
    if(destProcID == 29) return 573;
    if(destProcID == 38) return 574;
    if(destProcID == 46) return 575;
    if(destProcID == 60) return 576;
    if(destProcID == 64) return 577;
    if(destProcID == 107) return 578;
    if(destProcID == 114) return 579;
    if(destProcID == 120) return 580;
    if(destProcID == 130) return 581;
    if(destProcID == 2) return 582;
    if(destProcID == 25) return 583;
    if(destProcID == 23) return 584;
    if(destProcID == 14) return 585;
    if(destProcID == 6) return 586;
    if(destProcID == 125) return 587;
    if(destProcID == 121) return 588;
    if(destProcID == 78) return 589;
    if(destProcID == 71) return 590;
    if(destProcID == 65) return 591;
    if(destProcID == 55) return 592;
    if(destProcID == 50) return 593;
  end
  if (srcProcId == 27) begin
    if(destProcID == 28) return 594;
    if(destProcID == 30) return 595;
    if(destProcID == 39) return 596;
    if(destProcID == 47) return 597;
    if(destProcID == 61) return 598;
    if(destProcID == 65) return 599;
    if(destProcID == 108) return 600;
    if(destProcID == 115) return 601;
    if(destProcID == 121) return 602;
    if(destProcID == 131) return 603;
    if(destProcID == 3) return 604;
    if(destProcID == 26) return 605;
    if(destProcID == 24) return 606;
    if(destProcID == 15) return 607;
    if(destProcID == 7) return 608;
    if(destProcID == 126) return 609;
    if(destProcID == 122) return 610;
    if(destProcID == 79) return 611;
    if(destProcID == 72) return 612;
    if(destProcID == 66) return 613;
    if(destProcID == 56) return 614;
    if(destProcID == 51) return 615;
  end
  if (srcProcId == 28) begin
    if(destProcID == 29) return 616;
    if(destProcID == 31) return 617;
    if(destProcID == 40) return 618;
    if(destProcID == 48) return 619;
    if(destProcID == 62) return 620;
    if(destProcID == 66) return 621;
    if(destProcID == 109) return 622;
    if(destProcID == 116) return 623;
    if(destProcID == 122) return 624;
    if(destProcID == 132) return 625;
    if(destProcID == 4) return 626;
    if(destProcID == 27) return 627;
    if(destProcID == 25) return 628;
    if(destProcID == 16) return 629;
    if(destProcID == 8) return 630;
    if(destProcID == 127) return 631;
    if(destProcID == 123) return 632;
    if(destProcID == 80) return 633;
    if(destProcID == 73) return 634;
    if(destProcID == 67) return 635;
    if(destProcID == 57) return 636;
    if(destProcID == 52) return 637;
  end
  if (srcProcId == 29) begin
    if(destProcID == 30) return 638;
    if(destProcID == 32) return 639;
    if(destProcID == 41) return 640;
    if(destProcID == 49) return 641;
    if(destProcID == 63) return 642;
    if(destProcID == 67) return 643;
    if(destProcID == 110) return 644;
    if(destProcID == 117) return 645;
    if(destProcID == 123) return 646;
    if(destProcID == 0) return 647;
    if(destProcID == 5) return 648;
    if(destProcID == 28) return 649;
    if(destProcID == 26) return 650;
    if(destProcID == 17) return 651;
    if(destProcID == 9) return 652;
    if(destProcID == 128) return 653;
    if(destProcID == 124) return 654;
    if(destProcID == 81) return 655;
    if(destProcID == 74) return 656;
    if(destProcID == 68) return 657;
    if(destProcID == 58) return 658;
    if(destProcID == 53) return 659;
  end
  if (srcProcId == 30) begin
    if(destProcID == 31) return 660;
    if(destProcID == 33) return 661;
    if(destProcID == 42) return 662;
    if(destProcID == 50) return 663;
    if(destProcID == 64) return 664;
    if(destProcID == 68) return 665;
    if(destProcID == 111) return 666;
    if(destProcID == 118) return 667;
    if(destProcID == 124) return 668;
    if(destProcID == 1) return 669;
    if(destProcID == 6) return 670;
    if(destProcID == 29) return 671;
    if(destProcID == 27) return 672;
    if(destProcID == 18) return 673;
    if(destProcID == 10) return 674;
    if(destProcID == 129) return 675;
    if(destProcID == 125) return 676;
    if(destProcID == 82) return 677;
    if(destProcID == 75) return 678;
    if(destProcID == 69) return 679;
    if(destProcID == 59) return 680;
    if(destProcID == 54) return 681;
  end
  if (srcProcId == 31) begin
    if(destProcID == 32) return 682;
    if(destProcID == 34) return 683;
    if(destProcID == 43) return 684;
    if(destProcID == 51) return 685;
    if(destProcID == 65) return 686;
    if(destProcID == 69) return 687;
    if(destProcID == 112) return 688;
    if(destProcID == 119) return 689;
    if(destProcID == 125) return 690;
    if(destProcID == 2) return 691;
    if(destProcID == 7) return 692;
    if(destProcID == 30) return 693;
    if(destProcID == 28) return 694;
    if(destProcID == 19) return 695;
    if(destProcID == 11) return 696;
    if(destProcID == 130) return 697;
    if(destProcID == 126) return 698;
    if(destProcID == 83) return 699;
    if(destProcID == 76) return 700;
    if(destProcID == 70) return 701;
    if(destProcID == 60) return 702;
    if(destProcID == 55) return 703;
  end
  if (srcProcId == 32) begin
    if(destProcID == 33) return 704;
    if(destProcID == 35) return 705;
    if(destProcID == 44) return 706;
    if(destProcID == 52) return 707;
    if(destProcID == 66) return 708;
    if(destProcID == 70) return 709;
    if(destProcID == 113) return 710;
    if(destProcID == 120) return 711;
    if(destProcID == 126) return 712;
    if(destProcID == 3) return 713;
    if(destProcID == 8) return 714;
    if(destProcID == 31) return 715;
    if(destProcID == 29) return 716;
    if(destProcID == 20) return 717;
    if(destProcID == 12) return 718;
    if(destProcID == 131) return 719;
    if(destProcID == 127) return 720;
    if(destProcID == 84) return 721;
    if(destProcID == 77) return 722;
    if(destProcID == 71) return 723;
    if(destProcID == 61) return 724;
    if(destProcID == 56) return 725;
  end
  if (srcProcId == 33) begin
    if(destProcID == 34) return 726;
    if(destProcID == 36) return 727;
    if(destProcID == 45) return 728;
    if(destProcID == 53) return 729;
    if(destProcID == 67) return 730;
    if(destProcID == 71) return 731;
    if(destProcID == 114) return 732;
    if(destProcID == 121) return 733;
    if(destProcID == 127) return 734;
    if(destProcID == 4) return 735;
    if(destProcID == 9) return 736;
    if(destProcID == 32) return 737;
    if(destProcID == 30) return 738;
    if(destProcID == 21) return 739;
    if(destProcID == 13) return 740;
    if(destProcID == 132) return 741;
    if(destProcID == 128) return 742;
    if(destProcID == 85) return 743;
    if(destProcID == 78) return 744;
    if(destProcID == 72) return 745;
    if(destProcID == 62) return 746;
    if(destProcID == 57) return 747;
  end
  if (srcProcId == 34) begin
    if(destProcID == 35) return 748;
    if(destProcID == 37) return 749;
    if(destProcID == 46) return 750;
    if(destProcID == 54) return 751;
    if(destProcID == 68) return 752;
    if(destProcID == 72) return 753;
    if(destProcID == 115) return 754;
    if(destProcID == 122) return 755;
    if(destProcID == 128) return 756;
    if(destProcID == 5) return 757;
    if(destProcID == 10) return 758;
    if(destProcID == 33) return 759;
    if(destProcID == 31) return 760;
    if(destProcID == 22) return 761;
    if(destProcID == 14) return 762;
    if(destProcID == 0) return 763;
    if(destProcID == 129) return 764;
    if(destProcID == 86) return 765;
    if(destProcID == 79) return 766;
    if(destProcID == 73) return 767;
    if(destProcID == 63) return 768;
    if(destProcID == 58) return 769;
  end
  if (srcProcId == 35) begin
    if(destProcID == 36) return 770;
    if(destProcID == 38) return 771;
    if(destProcID == 47) return 772;
    if(destProcID == 55) return 773;
    if(destProcID == 69) return 774;
    if(destProcID == 73) return 775;
    if(destProcID == 116) return 776;
    if(destProcID == 123) return 777;
    if(destProcID == 129) return 778;
    if(destProcID == 6) return 779;
    if(destProcID == 11) return 780;
    if(destProcID == 34) return 781;
    if(destProcID == 32) return 782;
    if(destProcID == 23) return 783;
    if(destProcID == 15) return 784;
    if(destProcID == 1) return 785;
    if(destProcID == 130) return 786;
    if(destProcID == 87) return 787;
    if(destProcID == 80) return 788;
    if(destProcID == 74) return 789;
    if(destProcID == 64) return 790;
    if(destProcID == 59) return 791;
  end
  if (srcProcId == 36) begin
    if(destProcID == 37) return 792;
    if(destProcID == 39) return 793;
    if(destProcID == 48) return 794;
    if(destProcID == 56) return 795;
    if(destProcID == 70) return 796;
    if(destProcID == 74) return 797;
    if(destProcID == 117) return 798;
    if(destProcID == 124) return 799;
    if(destProcID == 130) return 800;
    if(destProcID == 7) return 801;
    if(destProcID == 12) return 802;
    if(destProcID == 35) return 803;
    if(destProcID == 33) return 804;
    if(destProcID == 24) return 805;
    if(destProcID == 16) return 806;
    if(destProcID == 2) return 807;
    if(destProcID == 131) return 808;
    if(destProcID == 88) return 809;
    if(destProcID == 81) return 810;
    if(destProcID == 75) return 811;
    if(destProcID == 65) return 812;
    if(destProcID == 60) return 813;
  end
  if (srcProcId == 37) begin
    if(destProcID == 38) return 814;
    if(destProcID == 40) return 815;
    if(destProcID == 49) return 816;
    if(destProcID == 57) return 817;
    if(destProcID == 71) return 818;
    if(destProcID == 75) return 819;
    if(destProcID == 118) return 820;
    if(destProcID == 125) return 821;
    if(destProcID == 131) return 822;
    if(destProcID == 8) return 823;
    if(destProcID == 13) return 824;
    if(destProcID == 36) return 825;
    if(destProcID == 34) return 826;
    if(destProcID == 25) return 827;
    if(destProcID == 17) return 828;
    if(destProcID == 3) return 829;
    if(destProcID == 132) return 830;
    if(destProcID == 89) return 831;
    if(destProcID == 82) return 832;
    if(destProcID == 76) return 833;
    if(destProcID == 66) return 834;
    if(destProcID == 61) return 835;
  end
  if (srcProcId == 38) begin
    if(destProcID == 39) return 836;
    if(destProcID == 41) return 837;
    if(destProcID == 50) return 838;
    if(destProcID == 58) return 839;
    if(destProcID == 72) return 840;
    if(destProcID == 76) return 841;
    if(destProcID == 119) return 842;
    if(destProcID == 126) return 843;
    if(destProcID == 132) return 844;
    if(destProcID == 9) return 845;
    if(destProcID == 14) return 846;
    if(destProcID == 37) return 847;
    if(destProcID == 35) return 848;
    if(destProcID == 26) return 849;
    if(destProcID == 18) return 850;
    if(destProcID == 4) return 851;
    if(destProcID == 0) return 852;
    if(destProcID == 90) return 853;
    if(destProcID == 83) return 854;
    if(destProcID == 77) return 855;
    if(destProcID == 67) return 856;
    if(destProcID == 62) return 857;
  end
  if (srcProcId == 39) begin
    if(destProcID == 40) return 858;
    if(destProcID == 42) return 859;
    if(destProcID == 51) return 860;
    if(destProcID == 59) return 861;
    if(destProcID == 73) return 862;
    if(destProcID == 77) return 863;
    if(destProcID == 120) return 864;
    if(destProcID == 127) return 865;
    if(destProcID == 0) return 866;
    if(destProcID == 10) return 867;
    if(destProcID == 15) return 868;
    if(destProcID == 38) return 869;
    if(destProcID == 36) return 870;
    if(destProcID == 27) return 871;
    if(destProcID == 19) return 872;
    if(destProcID == 5) return 873;
    if(destProcID == 1) return 874;
    if(destProcID == 91) return 875;
    if(destProcID == 84) return 876;
    if(destProcID == 78) return 877;
    if(destProcID == 68) return 878;
    if(destProcID == 63) return 879;
  end
  if (srcProcId == 40) begin
    if(destProcID == 41) return 880;
    if(destProcID == 43) return 881;
    if(destProcID == 52) return 882;
    if(destProcID == 60) return 883;
    if(destProcID == 74) return 884;
    if(destProcID == 78) return 885;
    if(destProcID == 121) return 886;
    if(destProcID == 128) return 887;
    if(destProcID == 1) return 888;
    if(destProcID == 11) return 889;
    if(destProcID == 16) return 890;
    if(destProcID == 39) return 891;
    if(destProcID == 37) return 892;
    if(destProcID == 28) return 893;
    if(destProcID == 20) return 894;
    if(destProcID == 6) return 895;
    if(destProcID == 2) return 896;
    if(destProcID == 92) return 897;
    if(destProcID == 85) return 898;
    if(destProcID == 79) return 899;
    if(destProcID == 69) return 900;
    if(destProcID == 64) return 901;
  end
  if (srcProcId == 41) begin
    if(destProcID == 42) return 902;
    if(destProcID == 44) return 903;
    if(destProcID == 53) return 904;
    if(destProcID == 61) return 905;
    if(destProcID == 75) return 906;
    if(destProcID == 79) return 907;
    if(destProcID == 122) return 908;
    if(destProcID == 129) return 909;
    if(destProcID == 2) return 910;
    if(destProcID == 12) return 911;
    if(destProcID == 17) return 912;
    if(destProcID == 40) return 913;
    if(destProcID == 38) return 914;
    if(destProcID == 29) return 915;
    if(destProcID == 21) return 916;
    if(destProcID == 7) return 917;
    if(destProcID == 3) return 918;
    if(destProcID == 93) return 919;
    if(destProcID == 86) return 920;
    if(destProcID == 80) return 921;
    if(destProcID == 70) return 922;
    if(destProcID == 65) return 923;
  end
  if (srcProcId == 42) begin
    if(destProcID == 43) return 924;
    if(destProcID == 45) return 925;
    if(destProcID == 54) return 926;
    if(destProcID == 62) return 927;
    if(destProcID == 76) return 928;
    if(destProcID == 80) return 929;
    if(destProcID == 123) return 930;
    if(destProcID == 130) return 931;
    if(destProcID == 3) return 932;
    if(destProcID == 13) return 933;
    if(destProcID == 18) return 934;
    if(destProcID == 41) return 935;
    if(destProcID == 39) return 936;
    if(destProcID == 30) return 937;
    if(destProcID == 22) return 938;
    if(destProcID == 8) return 939;
    if(destProcID == 4) return 940;
    if(destProcID == 94) return 941;
    if(destProcID == 87) return 942;
    if(destProcID == 81) return 943;
    if(destProcID == 71) return 944;
    if(destProcID == 66) return 945;
  end
  if (srcProcId == 43) begin
    if(destProcID == 44) return 946;
    if(destProcID == 46) return 947;
    if(destProcID == 55) return 948;
    if(destProcID == 63) return 949;
    if(destProcID == 77) return 950;
    if(destProcID == 81) return 951;
    if(destProcID == 124) return 952;
    if(destProcID == 131) return 953;
    if(destProcID == 4) return 954;
    if(destProcID == 14) return 955;
    if(destProcID == 19) return 956;
    if(destProcID == 42) return 957;
    if(destProcID == 40) return 958;
    if(destProcID == 31) return 959;
    if(destProcID == 23) return 960;
    if(destProcID == 9) return 961;
    if(destProcID == 5) return 962;
    if(destProcID == 95) return 963;
    if(destProcID == 88) return 964;
    if(destProcID == 82) return 965;
    if(destProcID == 72) return 966;
    if(destProcID == 67) return 967;
  end
  if (srcProcId == 44) begin
    if(destProcID == 45) return 968;
    if(destProcID == 47) return 969;
    if(destProcID == 56) return 970;
    if(destProcID == 64) return 971;
    if(destProcID == 78) return 972;
    if(destProcID == 82) return 973;
    if(destProcID == 125) return 974;
    if(destProcID == 132) return 975;
    if(destProcID == 5) return 976;
    if(destProcID == 15) return 977;
    if(destProcID == 20) return 978;
    if(destProcID == 43) return 979;
    if(destProcID == 41) return 980;
    if(destProcID == 32) return 981;
    if(destProcID == 24) return 982;
    if(destProcID == 10) return 983;
    if(destProcID == 6) return 984;
    if(destProcID == 96) return 985;
    if(destProcID == 89) return 986;
    if(destProcID == 83) return 987;
    if(destProcID == 73) return 988;
    if(destProcID == 68) return 989;
  end
  if (srcProcId == 45) begin
    if(destProcID == 46) return 990;
    if(destProcID == 48) return 991;
    if(destProcID == 57) return 992;
    if(destProcID == 65) return 993;
    if(destProcID == 79) return 994;
    if(destProcID == 83) return 995;
    if(destProcID == 126) return 996;
    if(destProcID == 0) return 997;
    if(destProcID == 6) return 998;
    if(destProcID == 16) return 999;
    if(destProcID == 21) return 1000;
    if(destProcID == 44) return 1001;
    if(destProcID == 42) return 1002;
    if(destProcID == 33) return 1003;
    if(destProcID == 25) return 1004;
    if(destProcID == 11) return 1005;
    if(destProcID == 7) return 1006;
    if(destProcID == 97) return 1007;
    if(destProcID == 90) return 1008;
    if(destProcID == 84) return 1009;
    if(destProcID == 74) return 1010;
    if(destProcID == 69) return 1011;
  end
  if (srcProcId == 46) begin
    if(destProcID == 47) return 1012;
    if(destProcID == 49) return 1013;
    if(destProcID == 58) return 1014;
    if(destProcID == 66) return 1015;
    if(destProcID == 80) return 1016;
    if(destProcID == 84) return 1017;
    if(destProcID == 127) return 1018;
    if(destProcID == 1) return 1019;
    if(destProcID == 7) return 1020;
    if(destProcID == 17) return 1021;
    if(destProcID == 22) return 1022;
    if(destProcID == 45) return 1023;
    if(destProcID == 43) return 1024;
    if(destProcID == 34) return 1025;
    if(destProcID == 26) return 1026;
    if(destProcID == 12) return 1027;
    if(destProcID == 8) return 1028;
    if(destProcID == 98) return 1029;
    if(destProcID == 91) return 1030;
    if(destProcID == 85) return 1031;
    if(destProcID == 75) return 1032;
    if(destProcID == 70) return 1033;
  end
  if (srcProcId == 47) begin
    if(destProcID == 48) return 1034;
    if(destProcID == 50) return 1035;
    if(destProcID == 59) return 1036;
    if(destProcID == 67) return 1037;
    if(destProcID == 81) return 1038;
    if(destProcID == 85) return 1039;
    if(destProcID == 128) return 1040;
    if(destProcID == 2) return 1041;
    if(destProcID == 8) return 1042;
    if(destProcID == 18) return 1043;
    if(destProcID == 23) return 1044;
    if(destProcID == 46) return 1045;
    if(destProcID == 44) return 1046;
    if(destProcID == 35) return 1047;
    if(destProcID == 27) return 1048;
    if(destProcID == 13) return 1049;
    if(destProcID == 9) return 1050;
    if(destProcID == 99) return 1051;
    if(destProcID == 92) return 1052;
    if(destProcID == 86) return 1053;
    if(destProcID == 76) return 1054;
    if(destProcID == 71) return 1055;
  end
  if (srcProcId == 48) begin
    if(destProcID == 49) return 1056;
    if(destProcID == 51) return 1057;
    if(destProcID == 60) return 1058;
    if(destProcID == 68) return 1059;
    if(destProcID == 82) return 1060;
    if(destProcID == 86) return 1061;
    if(destProcID == 129) return 1062;
    if(destProcID == 3) return 1063;
    if(destProcID == 9) return 1064;
    if(destProcID == 19) return 1065;
    if(destProcID == 24) return 1066;
    if(destProcID == 47) return 1067;
    if(destProcID == 45) return 1068;
    if(destProcID == 36) return 1069;
    if(destProcID == 28) return 1070;
    if(destProcID == 14) return 1071;
    if(destProcID == 10) return 1072;
    if(destProcID == 100) return 1073;
    if(destProcID == 93) return 1074;
    if(destProcID == 87) return 1075;
    if(destProcID == 77) return 1076;
    if(destProcID == 72) return 1077;
  end
  if (srcProcId == 49) begin
    if(destProcID == 50) return 1078;
    if(destProcID == 52) return 1079;
    if(destProcID == 61) return 1080;
    if(destProcID == 69) return 1081;
    if(destProcID == 83) return 1082;
    if(destProcID == 87) return 1083;
    if(destProcID == 130) return 1084;
    if(destProcID == 4) return 1085;
    if(destProcID == 10) return 1086;
    if(destProcID == 20) return 1087;
    if(destProcID == 25) return 1088;
    if(destProcID == 48) return 1089;
    if(destProcID == 46) return 1090;
    if(destProcID == 37) return 1091;
    if(destProcID == 29) return 1092;
    if(destProcID == 15) return 1093;
    if(destProcID == 11) return 1094;
    if(destProcID == 101) return 1095;
    if(destProcID == 94) return 1096;
    if(destProcID == 88) return 1097;
    if(destProcID == 78) return 1098;
    if(destProcID == 73) return 1099;
  end
  if (srcProcId == 50) begin
    if(destProcID == 51) return 1100;
    if(destProcID == 53) return 1101;
    if(destProcID == 62) return 1102;
    if(destProcID == 70) return 1103;
    if(destProcID == 84) return 1104;
    if(destProcID == 88) return 1105;
    if(destProcID == 131) return 1106;
    if(destProcID == 5) return 1107;
    if(destProcID == 11) return 1108;
    if(destProcID == 21) return 1109;
    if(destProcID == 26) return 1110;
    if(destProcID == 49) return 1111;
    if(destProcID == 47) return 1112;
    if(destProcID == 38) return 1113;
    if(destProcID == 30) return 1114;
    if(destProcID == 16) return 1115;
    if(destProcID == 12) return 1116;
    if(destProcID == 102) return 1117;
    if(destProcID == 95) return 1118;
    if(destProcID == 89) return 1119;
    if(destProcID == 79) return 1120;
    if(destProcID == 74) return 1121;
  end
  if (srcProcId == 51) begin
    if(destProcID == 52) return 1122;
    if(destProcID == 54) return 1123;
    if(destProcID == 63) return 1124;
    if(destProcID == 71) return 1125;
    if(destProcID == 85) return 1126;
    if(destProcID == 89) return 1127;
    if(destProcID == 132) return 1128;
    if(destProcID == 6) return 1129;
    if(destProcID == 12) return 1130;
    if(destProcID == 22) return 1131;
    if(destProcID == 27) return 1132;
    if(destProcID == 50) return 1133;
    if(destProcID == 48) return 1134;
    if(destProcID == 39) return 1135;
    if(destProcID == 31) return 1136;
    if(destProcID == 17) return 1137;
    if(destProcID == 13) return 1138;
    if(destProcID == 103) return 1139;
    if(destProcID == 96) return 1140;
    if(destProcID == 90) return 1141;
    if(destProcID == 80) return 1142;
    if(destProcID == 75) return 1143;
  end
  if (srcProcId == 52) begin
    if(destProcID == 53) return 1144;
    if(destProcID == 55) return 1145;
    if(destProcID == 64) return 1146;
    if(destProcID == 72) return 1147;
    if(destProcID == 86) return 1148;
    if(destProcID == 90) return 1149;
    if(destProcID == 0) return 1150;
    if(destProcID == 7) return 1151;
    if(destProcID == 13) return 1152;
    if(destProcID == 23) return 1153;
    if(destProcID == 28) return 1154;
    if(destProcID == 51) return 1155;
    if(destProcID == 49) return 1156;
    if(destProcID == 40) return 1157;
    if(destProcID == 32) return 1158;
    if(destProcID == 18) return 1159;
    if(destProcID == 14) return 1160;
    if(destProcID == 104) return 1161;
    if(destProcID == 97) return 1162;
    if(destProcID == 91) return 1163;
    if(destProcID == 81) return 1164;
    if(destProcID == 76) return 1165;
  end
  if (srcProcId == 53) begin
    if(destProcID == 54) return 1166;
    if(destProcID == 56) return 1167;
    if(destProcID == 65) return 1168;
    if(destProcID == 73) return 1169;
    if(destProcID == 87) return 1170;
    if(destProcID == 91) return 1171;
    if(destProcID == 1) return 1172;
    if(destProcID == 8) return 1173;
    if(destProcID == 14) return 1174;
    if(destProcID == 24) return 1175;
    if(destProcID == 29) return 1176;
    if(destProcID == 52) return 1177;
    if(destProcID == 50) return 1178;
    if(destProcID == 41) return 1179;
    if(destProcID == 33) return 1180;
    if(destProcID == 19) return 1181;
    if(destProcID == 15) return 1182;
    if(destProcID == 105) return 1183;
    if(destProcID == 98) return 1184;
    if(destProcID == 92) return 1185;
    if(destProcID == 82) return 1186;
    if(destProcID == 77) return 1187;
  end
  if (srcProcId == 54) begin
    if(destProcID == 55) return 1188;
    if(destProcID == 57) return 1189;
    if(destProcID == 66) return 1190;
    if(destProcID == 74) return 1191;
    if(destProcID == 88) return 1192;
    if(destProcID == 92) return 1193;
    if(destProcID == 2) return 1194;
    if(destProcID == 9) return 1195;
    if(destProcID == 15) return 1196;
    if(destProcID == 25) return 1197;
    if(destProcID == 30) return 1198;
    if(destProcID == 53) return 1199;
    if(destProcID == 51) return 1200;
    if(destProcID == 42) return 1201;
    if(destProcID == 34) return 1202;
    if(destProcID == 20) return 1203;
    if(destProcID == 16) return 1204;
    if(destProcID == 106) return 1205;
    if(destProcID == 99) return 1206;
    if(destProcID == 93) return 1207;
    if(destProcID == 83) return 1208;
    if(destProcID == 78) return 1209;
  end
  if (srcProcId == 55) begin
    if(destProcID == 56) return 1210;
    if(destProcID == 58) return 1211;
    if(destProcID == 67) return 1212;
    if(destProcID == 75) return 1213;
    if(destProcID == 89) return 1214;
    if(destProcID == 93) return 1215;
    if(destProcID == 3) return 1216;
    if(destProcID == 10) return 1217;
    if(destProcID == 16) return 1218;
    if(destProcID == 26) return 1219;
    if(destProcID == 31) return 1220;
    if(destProcID == 54) return 1221;
    if(destProcID == 52) return 1222;
    if(destProcID == 43) return 1223;
    if(destProcID == 35) return 1224;
    if(destProcID == 21) return 1225;
    if(destProcID == 17) return 1226;
    if(destProcID == 107) return 1227;
    if(destProcID == 100) return 1228;
    if(destProcID == 94) return 1229;
    if(destProcID == 84) return 1230;
    if(destProcID == 79) return 1231;
  end
  if (srcProcId == 56) begin
    if(destProcID == 57) return 1232;
    if(destProcID == 59) return 1233;
    if(destProcID == 68) return 1234;
    if(destProcID == 76) return 1235;
    if(destProcID == 90) return 1236;
    if(destProcID == 94) return 1237;
    if(destProcID == 4) return 1238;
    if(destProcID == 11) return 1239;
    if(destProcID == 17) return 1240;
    if(destProcID == 27) return 1241;
    if(destProcID == 32) return 1242;
    if(destProcID == 55) return 1243;
    if(destProcID == 53) return 1244;
    if(destProcID == 44) return 1245;
    if(destProcID == 36) return 1246;
    if(destProcID == 22) return 1247;
    if(destProcID == 18) return 1248;
    if(destProcID == 108) return 1249;
    if(destProcID == 101) return 1250;
    if(destProcID == 95) return 1251;
    if(destProcID == 85) return 1252;
    if(destProcID == 80) return 1253;
  end
  if (srcProcId == 57) begin
    if(destProcID == 58) return 1254;
    if(destProcID == 60) return 1255;
    if(destProcID == 69) return 1256;
    if(destProcID == 77) return 1257;
    if(destProcID == 91) return 1258;
    if(destProcID == 95) return 1259;
    if(destProcID == 5) return 1260;
    if(destProcID == 12) return 1261;
    if(destProcID == 18) return 1262;
    if(destProcID == 28) return 1263;
    if(destProcID == 33) return 1264;
    if(destProcID == 56) return 1265;
    if(destProcID == 54) return 1266;
    if(destProcID == 45) return 1267;
    if(destProcID == 37) return 1268;
    if(destProcID == 23) return 1269;
    if(destProcID == 19) return 1270;
    if(destProcID == 109) return 1271;
    if(destProcID == 102) return 1272;
    if(destProcID == 96) return 1273;
    if(destProcID == 86) return 1274;
    if(destProcID == 81) return 1275;
  end
  if (srcProcId == 58) begin
    if(destProcID == 59) return 1276;
    if(destProcID == 61) return 1277;
    if(destProcID == 70) return 1278;
    if(destProcID == 78) return 1279;
    if(destProcID == 92) return 1280;
    if(destProcID == 96) return 1281;
    if(destProcID == 6) return 1282;
    if(destProcID == 13) return 1283;
    if(destProcID == 19) return 1284;
    if(destProcID == 29) return 1285;
    if(destProcID == 34) return 1286;
    if(destProcID == 57) return 1287;
    if(destProcID == 55) return 1288;
    if(destProcID == 46) return 1289;
    if(destProcID == 38) return 1290;
    if(destProcID == 24) return 1291;
    if(destProcID == 20) return 1292;
    if(destProcID == 110) return 1293;
    if(destProcID == 103) return 1294;
    if(destProcID == 97) return 1295;
    if(destProcID == 87) return 1296;
    if(destProcID == 82) return 1297;
  end
  if (srcProcId == 59) begin
    if(destProcID == 60) return 1298;
    if(destProcID == 62) return 1299;
    if(destProcID == 71) return 1300;
    if(destProcID == 79) return 1301;
    if(destProcID == 93) return 1302;
    if(destProcID == 97) return 1303;
    if(destProcID == 7) return 1304;
    if(destProcID == 14) return 1305;
    if(destProcID == 20) return 1306;
    if(destProcID == 30) return 1307;
    if(destProcID == 35) return 1308;
    if(destProcID == 58) return 1309;
    if(destProcID == 56) return 1310;
    if(destProcID == 47) return 1311;
    if(destProcID == 39) return 1312;
    if(destProcID == 25) return 1313;
    if(destProcID == 21) return 1314;
    if(destProcID == 111) return 1315;
    if(destProcID == 104) return 1316;
    if(destProcID == 98) return 1317;
    if(destProcID == 88) return 1318;
    if(destProcID == 83) return 1319;
  end
  if (srcProcId == 60) begin
    if(destProcID == 61) return 1320;
    if(destProcID == 63) return 1321;
    if(destProcID == 72) return 1322;
    if(destProcID == 80) return 1323;
    if(destProcID == 94) return 1324;
    if(destProcID == 98) return 1325;
    if(destProcID == 8) return 1326;
    if(destProcID == 15) return 1327;
    if(destProcID == 21) return 1328;
    if(destProcID == 31) return 1329;
    if(destProcID == 36) return 1330;
    if(destProcID == 59) return 1331;
    if(destProcID == 57) return 1332;
    if(destProcID == 48) return 1333;
    if(destProcID == 40) return 1334;
    if(destProcID == 26) return 1335;
    if(destProcID == 22) return 1336;
    if(destProcID == 112) return 1337;
    if(destProcID == 105) return 1338;
    if(destProcID == 99) return 1339;
    if(destProcID == 89) return 1340;
    if(destProcID == 84) return 1341;
  end
  if (srcProcId == 61) begin
    if(destProcID == 62) return 1342;
    if(destProcID == 64) return 1343;
    if(destProcID == 73) return 1344;
    if(destProcID == 81) return 1345;
    if(destProcID == 95) return 1346;
    if(destProcID == 99) return 1347;
    if(destProcID == 9) return 1348;
    if(destProcID == 16) return 1349;
    if(destProcID == 22) return 1350;
    if(destProcID == 32) return 1351;
    if(destProcID == 37) return 1352;
    if(destProcID == 60) return 1353;
    if(destProcID == 58) return 1354;
    if(destProcID == 49) return 1355;
    if(destProcID == 41) return 1356;
    if(destProcID == 27) return 1357;
    if(destProcID == 23) return 1358;
    if(destProcID == 113) return 1359;
    if(destProcID == 106) return 1360;
    if(destProcID == 100) return 1361;
    if(destProcID == 90) return 1362;
    if(destProcID == 85) return 1363;
  end
  if (srcProcId == 62) begin
    if(destProcID == 63) return 1364;
    if(destProcID == 65) return 1365;
    if(destProcID == 74) return 1366;
    if(destProcID == 82) return 1367;
    if(destProcID == 96) return 1368;
    if(destProcID == 100) return 1369;
    if(destProcID == 10) return 1370;
    if(destProcID == 17) return 1371;
    if(destProcID == 23) return 1372;
    if(destProcID == 33) return 1373;
    if(destProcID == 38) return 1374;
    if(destProcID == 61) return 1375;
    if(destProcID == 59) return 1376;
    if(destProcID == 50) return 1377;
    if(destProcID == 42) return 1378;
    if(destProcID == 28) return 1379;
    if(destProcID == 24) return 1380;
    if(destProcID == 114) return 1381;
    if(destProcID == 107) return 1382;
    if(destProcID == 101) return 1383;
    if(destProcID == 91) return 1384;
    if(destProcID == 86) return 1385;
  end
  if (srcProcId == 63) begin
    if(destProcID == 64) return 1386;
    if(destProcID == 66) return 1387;
    if(destProcID == 75) return 1388;
    if(destProcID == 83) return 1389;
    if(destProcID == 97) return 1390;
    if(destProcID == 101) return 1391;
    if(destProcID == 11) return 1392;
    if(destProcID == 18) return 1393;
    if(destProcID == 24) return 1394;
    if(destProcID == 34) return 1395;
    if(destProcID == 39) return 1396;
    if(destProcID == 62) return 1397;
    if(destProcID == 60) return 1398;
    if(destProcID == 51) return 1399;
    if(destProcID == 43) return 1400;
    if(destProcID == 29) return 1401;
    if(destProcID == 25) return 1402;
    if(destProcID == 115) return 1403;
    if(destProcID == 108) return 1404;
    if(destProcID == 102) return 1405;
    if(destProcID == 92) return 1406;
    if(destProcID == 87) return 1407;
  end
  if (srcProcId == 64) begin
    if(destProcID == 65) return 1408;
    if(destProcID == 67) return 1409;
    if(destProcID == 76) return 1410;
    if(destProcID == 84) return 1411;
    if(destProcID == 98) return 1412;
    if(destProcID == 102) return 1413;
    if(destProcID == 12) return 1414;
    if(destProcID == 19) return 1415;
    if(destProcID == 25) return 1416;
    if(destProcID == 35) return 1417;
    if(destProcID == 40) return 1418;
    if(destProcID == 63) return 1419;
    if(destProcID == 61) return 1420;
    if(destProcID == 52) return 1421;
    if(destProcID == 44) return 1422;
    if(destProcID == 30) return 1423;
    if(destProcID == 26) return 1424;
    if(destProcID == 116) return 1425;
    if(destProcID == 109) return 1426;
    if(destProcID == 103) return 1427;
    if(destProcID == 93) return 1428;
    if(destProcID == 88) return 1429;
  end
  if (srcProcId == 65) begin
    if(destProcID == 66) return 1430;
    if(destProcID == 68) return 1431;
    if(destProcID == 77) return 1432;
    if(destProcID == 85) return 1433;
    if(destProcID == 99) return 1434;
    if(destProcID == 103) return 1435;
    if(destProcID == 13) return 1436;
    if(destProcID == 20) return 1437;
    if(destProcID == 26) return 1438;
    if(destProcID == 36) return 1439;
    if(destProcID == 41) return 1440;
    if(destProcID == 64) return 1441;
    if(destProcID == 62) return 1442;
    if(destProcID == 53) return 1443;
    if(destProcID == 45) return 1444;
    if(destProcID == 31) return 1445;
    if(destProcID == 27) return 1446;
    if(destProcID == 117) return 1447;
    if(destProcID == 110) return 1448;
    if(destProcID == 104) return 1449;
    if(destProcID == 94) return 1450;
    if(destProcID == 89) return 1451;
  end
  if (srcProcId == 66) begin
    if(destProcID == 67) return 1452;
    if(destProcID == 69) return 1453;
    if(destProcID == 78) return 1454;
    if(destProcID == 86) return 1455;
    if(destProcID == 100) return 1456;
    if(destProcID == 104) return 1457;
    if(destProcID == 14) return 1458;
    if(destProcID == 21) return 1459;
    if(destProcID == 27) return 1460;
    if(destProcID == 37) return 1461;
    if(destProcID == 42) return 1462;
    if(destProcID == 65) return 1463;
    if(destProcID == 63) return 1464;
    if(destProcID == 54) return 1465;
    if(destProcID == 46) return 1466;
    if(destProcID == 32) return 1467;
    if(destProcID == 28) return 1468;
    if(destProcID == 118) return 1469;
    if(destProcID == 111) return 1470;
    if(destProcID == 105) return 1471;
    if(destProcID == 95) return 1472;
    if(destProcID == 90) return 1473;
  end
  if (srcProcId == 67) begin
    if(destProcID == 68) return 1474;
    if(destProcID == 70) return 1475;
    if(destProcID == 79) return 1476;
    if(destProcID == 87) return 1477;
    if(destProcID == 101) return 1478;
    if(destProcID == 105) return 1479;
    if(destProcID == 15) return 1480;
    if(destProcID == 22) return 1481;
    if(destProcID == 28) return 1482;
    if(destProcID == 38) return 1483;
    if(destProcID == 43) return 1484;
    if(destProcID == 66) return 1485;
    if(destProcID == 64) return 1486;
    if(destProcID == 55) return 1487;
    if(destProcID == 47) return 1488;
    if(destProcID == 33) return 1489;
    if(destProcID == 29) return 1490;
    if(destProcID == 119) return 1491;
    if(destProcID == 112) return 1492;
    if(destProcID == 106) return 1493;
    if(destProcID == 96) return 1494;
    if(destProcID == 91) return 1495;
  end
  if (srcProcId == 68) begin
    if(destProcID == 69) return 1496;
    if(destProcID == 71) return 1497;
    if(destProcID == 80) return 1498;
    if(destProcID == 88) return 1499;
    if(destProcID == 102) return 1500;
    if(destProcID == 106) return 1501;
    if(destProcID == 16) return 1502;
    if(destProcID == 23) return 1503;
    if(destProcID == 29) return 1504;
    if(destProcID == 39) return 1505;
    if(destProcID == 44) return 1506;
    if(destProcID == 67) return 1507;
    if(destProcID == 65) return 1508;
    if(destProcID == 56) return 1509;
    if(destProcID == 48) return 1510;
    if(destProcID == 34) return 1511;
    if(destProcID == 30) return 1512;
    if(destProcID == 120) return 1513;
    if(destProcID == 113) return 1514;
    if(destProcID == 107) return 1515;
    if(destProcID == 97) return 1516;
    if(destProcID == 92) return 1517;
  end
  if (srcProcId == 69) begin
    if(destProcID == 70) return 1518;
    if(destProcID == 72) return 1519;
    if(destProcID == 81) return 1520;
    if(destProcID == 89) return 1521;
    if(destProcID == 103) return 1522;
    if(destProcID == 107) return 1523;
    if(destProcID == 17) return 1524;
    if(destProcID == 24) return 1525;
    if(destProcID == 30) return 1526;
    if(destProcID == 40) return 1527;
    if(destProcID == 45) return 1528;
    if(destProcID == 68) return 1529;
    if(destProcID == 66) return 1530;
    if(destProcID == 57) return 1531;
    if(destProcID == 49) return 1532;
    if(destProcID == 35) return 1533;
    if(destProcID == 31) return 1534;
    if(destProcID == 121) return 1535;
    if(destProcID == 114) return 1536;
    if(destProcID == 108) return 1537;
    if(destProcID == 98) return 1538;
    if(destProcID == 93) return 1539;
  end
  if (srcProcId == 70) begin
    if(destProcID == 71) return 1540;
    if(destProcID == 73) return 1541;
    if(destProcID == 82) return 1542;
    if(destProcID == 90) return 1543;
    if(destProcID == 104) return 1544;
    if(destProcID == 108) return 1545;
    if(destProcID == 18) return 1546;
    if(destProcID == 25) return 1547;
    if(destProcID == 31) return 1548;
    if(destProcID == 41) return 1549;
    if(destProcID == 46) return 1550;
    if(destProcID == 69) return 1551;
    if(destProcID == 67) return 1552;
    if(destProcID == 58) return 1553;
    if(destProcID == 50) return 1554;
    if(destProcID == 36) return 1555;
    if(destProcID == 32) return 1556;
    if(destProcID == 122) return 1557;
    if(destProcID == 115) return 1558;
    if(destProcID == 109) return 1559;
    if(destProcID == 99) return 1560;
    if(destProcID == 94) return 1561;
  end
  if (srcProcId == 71) begin
    if(destProcID == 72) return 1562;
    if(destProcID == 74) return 1563;
    if(destProcID == 83) return 1564;
    if(destProcID == 91) return 1565;
    if(destProcID == 105) return 1566;
    if(destProcID == 109) return 1567;
    if(destProcID == 19) return 1568;
    if(destProcID == 26) return 1569;
    if(destProcID == 32) return 1570;
    if(destProcID == 42) return 1571;
    if(destProcID == 47) return 1572;
    if(destProcID == 70) return 1573;
    if(destProcID == 68) return 1574;
    if(destProcID == 59) return 1575;
    if(destProcID == 51) return 1576;
    if(destProcID == 37) return 1577;
    if(destProcID == 33) return 1578;
    if(destProcID == 123) return 1579;
    if(destProcID == 116) return 1580;
    if(destProcID == 110) return 1581;
    if(destProcID == 100) return 1582;
    if(destProcID == 95) return 1583;
  end
  if (srcProcId == 72) begin
    if(destProcID == 73) return 1584;
    if(destProcID == 75) return 1585;
    if(destProcID == 84) return 1586;
    if(destProcID == 92) return 1587;
    if(destProcID == 106) return 1588;
    if(destProcID == 110) return 1589;
    if(destProcID == 20) return 1590;
    if(destProcID == 27) return 1591;
    if(destProcID == 33) return 1592;
    if(destProcID == 43) return 1593;
    if(destProcID == 48) return 1594;
    if(destProcID == 71) return 1595;
    if(destProcID == 69) return 1596;
    if(destProcID == 60) return 1597;
    if(destProcID == 52) return 1598;
    if(destProcID == 38) return 1599;
    if(destProcID == 34) return 1600;
    if(destProcID == 124) return 1601;
    if(destProcID == 117) return 1602;
    if(destProcID == 111) return 1603;
    if(destProcID == 101) return 1604;
    if(destProcID == 96) return 1605;
  end
  if (srcProcId == 73) begin
    if(destProcID == 74) return 1606;
    if(destProcID == 76) return 1607;
    if(destProcID == 85) return 1608;
    if(destProcID == 93) return 1609;
    if(destProcID == 107) return 1610;
    if(destProcID == 111) return 1611;
    if(destProcID == 21) return 1612;
    if(destProcID == 28) return 1613;
    if(destProcID == 34) return 1614;
    if(destProcID == 44) return 1615;
    if(destProcID == 49) return 1616;
    if(destProcID == 72) return 1617;
    if(destProcID == 70) return 1618;
    if(destProcID == 61) return 1619;
    if(destProcID == 53) return 1620;
    if(destProcID == 39) return 1621;
    if(destProcID == 35) return 1622;
    if(destProcID == 125) return 1623;
    if(destProcID == 118) return 1624;
    if(destProcID == 112) return 1625;
    if(destProcID == 102) return 1626;
    if(destProcID == 97) return 1627;
  end
  if (srcProcId == 74) begin
    if(destProcID == 75) return 1628;
    if(destProcID == 77) return 1629;
    if(destProcID == 86) return 1630;
    if(destProcID == 94) return 1631;
    if(destProcID == 108) return 1632;
    if(destProcID == 112) return 1633;
    if(destProcID == 22) return 1634;
    if(destProcID == 29) return 1635;
    if(destProcID == 35) return 1636;
    if(destProcID == 45) return 1637;
    if(destProcID == 50) return 1638;
    if(destProcID == 73) return 1639;
    if(destProcID == 71) return 1640;
    if(destProcID == 62) return 1641;
    if(destProcID == 54) return 1642;
    if(destProcID == 40) return 1643;
    if(destProcID == 36) return 1644;
    if(destProcID == 126) return 1645;
    if(destProcID == 119) return 1646;
    if(destProcID == 113) return 1647;
    if(destProcID == 103) return 1648;
    if(destProcID == 98) return 1649;
  end
  if (srcProcId == 75) begin
    if(destProcID == 76) return 1650;
    if(destProcID == 78) return 1651;
    if(destProcID == 87) return 1652;
    if(destProcID == 95) return 1653;
    if(destProcID == 109) return 1654;
    if(destProcID == 113) return 1655;
    if(destProcID == 23) return 1656;
    if(destProcID == 30) return 1657;
    if(destProcID == 36) return 1658;
    if(destProcID == 46) return 1659;
    if(destProcID == 51) return 1660;
    if(destProcID == 74) return 1661;
    if(destProcID == 72) return 1662;
    if(destProcID == 63) return 1663;
    if(destProcID == 55) return 1664;
    if(destProcID == 41) return 1665;
    if(destProcID == 37) return 1666;
    if(destProcID == 127) return 1667;
    if(destProcID == 120) return 1668;
    if(destProcID == 114) return 1669;
    if(destProcID == 104) return 1670;
    if(destProcID == 99) return 1671;
  end
  if (srcProcId == 76) begin
    if(destProcID == 77) return 1672;
    if(destProcID == 79) return 1673;
    if(destProcID == 88) return 1674;
    if(destProcID == 96) return 1675;
    if(destProcID == 110) return 1676;
    if(destProcID == 114) return 1677;
    if(destProcID == 24) return 1678;
    if(destProcID == 31) return 1679;
    if(destProcID == 37) return 1680;
    if(destProcID == 47) return 1681;
    if(destProcID == 52) return 1682;
    if(destProcID == 75) return 1683;
    if(destProcID == 73) return 1684;
    if(destProcID == 64) return 1685;
    if(destProcID == 56) return 1686;
    if(destProcID == 42) return 1687;
    if(destProcID == 38) return 1688;
    if(destProcID == 128) return 1689;
    if(destProcID == 121) return 1690;
    if(destProcID == 115) return 1691;
    if(destProcID == 105) return 1692;
    if(destProcID == 100) return 1693;
  end
  if (srcProcId == 77) begin
    if(destProcID == 78) return 1694;
    if(destProcID == 80) return 1695;
    if(destProcID == 89) return 1696;
    if(destProcID == 97) return 1697;
    if(destProcID == 111) return 1698;
    if(destProcID == 115) return 1699;
    if(destProcID == 25) return 1700;
    if(destProcID == 32) return 1701;
    if(destProcID == 38) return 1702;
    if(destProcID == 48) return 1703;
    if(destProcID == 53) return 1704;
    if(destProcID == 76) return 1705;
    if(destProcID == 74) return 1706;
    if(destProcID == 65) return 1707;
    if(destProcID == 57) return 1708;
    if(destProcID == 43) return 1709;
    if(destProcID == 39) return 1710;
    if(destProcID == 129) return 1711;
    if(destProcID == 122) return 1712;
    if(destProcID == 116) return 1713;
    if(destProcID == 106) return 1714;
    if(destProcID == 101) return 1715;
  end
  if (srcProcId == 78) begin
    if(destProcID == 79) return 1716;
    if(destProcID == 81) return 1717;
    if(destProcID == 90) return 1718;
    if(destProcID == 98) return 1719;
    if(destProcID == 112) return 1720;
    if(destProcID == 116) return 1721;
    if(destProcID == 26) return 1722;
    if(destProcID == 33) return 1723;
    if(destProcID == 39) return 1724;
    if(destProcID == 49) return 1725;
    if(destProcID == 54) return 1726;
    if(destProcID == 77) return 1727;
    if(destProcID == 75) return 1728;
    if(destProcID == 66) return 1729;
    if(destProcID == 58) return 1730;
    if(destProcID == 44) return 1731;
    if(destProcID == 40) return 1732;
    if(destProcID == 130) return 1733;
    if(destProcID == 123) return 1734;
    if(destProcID == 117) return 1735;
    if(destProcID == 107) return 1736;
    if(destProcID == 102) return 1737;
  end
  if (srcProcId == 79) begin
    if(destProcID == 80) return 1738;
    if(destProcID == 82) return 1739;
    if(destProcID == 91) return 1740;
    if(destProcID == 99) return 1741;
    if(destProcID == 113) return 1742;
    if(destProcID == 117) return 1743;
    if(destProcID == 27) return 1744;
    if(destProcID == 34) return 1745;
    if(destProcID == 40) return 1746;
    if(destProcID == 50) return 1747;
    if(destProcID == 55) return 1748;
    if(destProcID == 78) return 1749;
    if(destProcID == 76) return 1750;
    if(destProcID == 67) return 1751;
    if(destProcID == 59) return 1752;
    if(destProcID == 45) return 1753;
    if(destProcID == 41) return 1754;
    if(destProcID == 131) return 1755;
    if(destProcID == 124) return 1756;
    if(destProcID == 118) return 1757;
    if(destProcID == 108) return 1758;
    if(destProcID == 103) return 1759;
  end
  if (srcProcId == 80) begin
    if(destProcID == 81) return 1760;
    if(destProcID == 83) return 1761;
    if(destProcID == 92) return 1762;
    if(destProcID == 100) return 1763;
    if(destProcID == 114) return 1764;
    if(destProcID == 118) return 1765;
    if(destProcID == 28) return 1766;
    if(destProcID == 35) return 1767;
    if(destProcID == 41) return 1768;
    if(destProcID == 51) return 1769;
    if(destProcID == 56) return 1770;
    if(destProcID == 79) return 1771;
    if(destProcID == 77) return 1772;
    if(destProcID == 68) return 1773;
    if(destProcID == 60) return 1774;
    if(destProcID == 46) return 1775;
    if(destProcID == 42) return 1776;
    if(destProcID == 132) return 1777;
    if(destProcID == 125) return 1778;
    if(destProcID == 119) return 1779;
    if(destProcID == 109) return 1780;
    if(destProcID == 104) return 1781;
  end
  if (srcProcId == 81) begin
    if(destProcID == 82) return 1782;
    if(destProcID == 84) return 1783;
    if(destProcID == 93) return 1784;
    if(destProcID == 101) return 1785;
    if(destProcID == 115) return 1786;
    if(destProcID == 119) return 1787;
    if(destProcID == 29) return 1788;
    if(destProcID == 36) return 1789;
    if(destProcID == 42) return 1790;
    if(destProcID == 52) return 1791;
    if(destProcID == 57) return 1792;
    if(destProcID == 80) return 1793;
    if(destProcID == 78) return 1794;
    if(destProcID == 69) return 1795;
    if(destProcID == 61) return 1796;
    if(destProcID == 47) return 1797;
    if(destProcID == 43) return 1798;
    if(destProcID == 0) return 1799;
    if(destProcID == 126) return 1800;
    if(destProcID == 120) return 1801;
    if(destProcID == 110) return 1802;
    if(destProcID == 105) return 1803;
  end
  if (srcProcId == 82) begin
    if(destProcID == 83) return 1804;
    if(destProcID == 85) return 1805;
    if(destProcID == 94) return 1806;
    if(destProcID == 102) return 1807;
    if(destProcID == 116) return 1808;
    if(destProcID == 120) return 1809;
    if(destProcID == 30) return 1810;
    if(destProcID == 37) return 1811;
    if(destProcID == 43) return 1812;
    if(destProcID == 53) return 1813;
    if(destProcID == 58) return 1814;
    if(destProcID == 81) return 1815;
    if(destProcID == 79) return 1816;
    if(destProcID == 70) return 1817;
    if(destProcID == 62) return 1818;
    if(destProcID == 48) return 1819;
    if(destProcID == 44) return 1820;
    if(destProcID == 1) return 1821;
    if(destProcID == 127) return 1822;
    if(destProcID == 121) return 1823;
    if(destProcID == 111) return 1824;
    if(destProcID == 106) return 1825;
  end
  if (srcProcId == 83) begin
    if(destProcID == 84) return 1826;
    if(destProcID == 86) return 1827;
    if(destProcID == 95) return 1828;
    if(destProcID == 103) return 1829;
    if(destProcID == 117) return 1830;
    if(destProcID == 121) return 1831;
    if(destProcID == 31) return 1832;
    if(destProcID == 38) return 1833;
    if(destProcID == 44) return 1834;
    if(destProcID == 54) return 1835;
    if(destProcID == 59) return 1836;
    if(destProcID == 82) return 1837;
    if(destProcID == 80) return 1838;
    if(destProcID == 71) return 1839;
    if(destProcID == 63) return 1840;
    if(destProcID == 49) return 1841;
    if(destProcID == 45) return 1842;
    if(destProcID == 2) return 1843;
    if(destProcID == 128) return 1844;
    if(destProcID == 122) return 1845;
    if(destProcID == 112) return 1846;
    if(destProcID == 107) return 1847;
  end
  if (srcProcId == 84) begin
    if(destProcID == 85) return 1848;
    if(destProcID == 87) return 1849;
    if(destProcID == 96) return 1850;
    if(destProcID == 104) return 1851;
    if(destProcID == 118) return 1852;
    if(destProcID == 122) return 1853;
    if(destProcID == 32) return 1854;
    if(destProcID == 39) return 1855;
    if(destProcID == 45) return 1856;
    if(destProcID == 55) return 1857;
    if(destProcID == 60) return 1858;
    if(destProcID == 83) return 1859;
    if(destProcID == 81) return 1860;
    if(destProcID == 72) return 1861;
    if(destProcID == 64) return 1862;
    if(destProcID == 50) return 1863;
    if(destProcID == 46) return 1864;
    if(destProcID == 3) return 1865;
    if(destProcID == 129) return 1866;
    if(destProcID == 123) return 1867;
    if(destProcID == 113) return 1868;
    if(destProcID == 108) return 1869;
  end
  if (srcProcId == 85) begin
    if(destProcID == 86) return 1870;
    if(destProcID == 88) return 1871;
    if(destProcID == 97) return 1872;
    if(destProcID == 105) return 1873;
    if(destProcID == 119) return 1874;
    if(destProcID == 123) return 1875;
    if(destProcID == 33) return 1876;
    if(destProcID == 40) return 1877;
    if(destProcID == 46) return 1878;
    if(destProcID == 56) return 1879;
    if(destProcID == 61) return 1880;
    if(destProcID == 84) return 1881;
    if(destProcID == 82) return 1882;
    if(destProcID == 73) return 1883;
    if(destProcID == 65) return 1884;
    if(destProcID == 51) return 1885;
    if(destProcID == 47) return 1886;
    if(destProcID == 4) return 1887;
    if(destProcID == 130) return 1888;
    if(destProcID == 124) return 1889;
    if(destProcID == 114) return 1890;
    if(destProcID == 109) return 1891;
  end
  if (srcProcId == 86) begin
    if(destProcID == 87) return 1892;
    if(destProcID == 89) return 1893;
    if(destProcID == 98) return 1894;
    if(destProcID == 106) return 1895;
    if(destProcID == 120) return 1896;
    if(destProcID == 124) return 1897;
    if(destProcID == 34) return 1898;
    if(destProcID == 41) return 1899;
    if(destProcID == 47) return 1900;
    if(destProcID == 57) return 1901;
    if(destProcID == 62) return 1902;
    if(destProcID == 85) return 1903;
    if(destProcID == 83) return 1904;
    if(destProcID == 74) return 1905;
    if(destProcID == 66) return 1906;
    if(destProcID == 52) return 1907;
    if(destProcID == 48) return 1908;
    if(destProcID == 5) return 1909;
    if(destProcID == 131) return 1910;
    if(destProcID == 125) return 1911;
    if(destProcID == 115) return 1912;
    if(destProcID == 110) return 1913;
  end
  if (srcProcId == 87) begin
    if(destProcID == 88) return 1914;
    if(destProcID == 90) return 1915;
    if(destProcID == 99) return 1916;
    if(destProcID == 107) return 1917;
    if(destProcID == 121) return 1918;
    if(destProcID == 125) return 1919;
    if(destProcID == 35) return 1920;
    if(destProcID == 42) return 1921;
    if(destProcID == 48) return 1922;
    if(destProcID == 58) return 1923;
    if(destProcID == 63) return 1924;
    if(destProcID == 86) return 1925;
    if(destProcID == 84) return 1926;
    if(destProcID == 75) return 1927;
    if(destProcID == 67) return 1928;
    if(destProcID == 53) return 1929;
    if(destProcID == 49) return 1930;
    if(destProcID == 6) return 1931;
    if(destProcID == 132) return 1932;
    if(destProcID == 126) return 1933;
    if(destProcID == 116) return 1934;
    if(destProcID == 111) return 1935;
  end
  if (srcProcId == 88) begin
    if(destProcID == 89) return 1936;
    if(destProcID == 91) return 1937;
    if(destProcID == 100) return 1938;
    if(destProcID == 108) return 1939;
    if(destProcID == 122) return 1940;
    if(destProcID == 126) return 1941;
    if(destProcID == 36) return 1942;
    if(destProcID == 43) return 1943;
    if(destProcID == 49) return 1944;
    if(destProcID == 59) return 1945;
    if(destProcID == 64) return 1946;
    if(destProcID == 87) return 1947;
    if(destProcID == 85) return 1948;
    if(destProcID == 76) return 1949;
    if(destProcID == 68) return 1950;
    if(destProcID == 54) return 1951;
    if(destProcID == 50) return 1952;
    if(destProcID == 7) return 1953;
    if(destProcID == 0) return 1954;
    if(destProcID == 127) return 1955;
    if(destProcID == 117) return 1956;
    if(destProcID == 112) return 1957;
  end
  if (srcProcId == 89) begin
    if(destProcID == 90) return 1958;
    if(destProcID == 92) return 1959;
    if(destProcID == 101) return 1960;
    if(destProcID == 109) return 1961;
    if(destProcID == 123) return 1962;
    if(destProcID == 127) return 1963;
    if(destProcID == 37) return 1964;
    if(destProcID == 44) return 1965;
    if(destProcID == 50) return 1966;
    if(destProcID == 60) return 1967;
    if(destProcID == 65) return 1968;
    if(destProcID == 88) return 1969;
    if(destProcID == 86) return 1970;
    if(destProcID == 77) return 1971;
    if(destProcID == 69) return 1972;
    if(destProcID == 55) return 1973;
    if(destProcID == 51) return 1974;
    if(destProcID == 8) return 1975;
    if(destProcID == 1) return 1976;
    if(destProcID == 128) return 1977;
    if(destProcID == 118) return 1978;
    if(destProcID == 113) return 1979;
  end
  if (srcProcId == 90) begin
    if(destProcID == 91) return 1980;
    if(destProcID == 93) return 1981;
    if(destProcID == 102) return 1982;
    if(destProcID == 110) return 1983;
    if(destProcID == 124) return 1984;
    if(destProcID == 128) return 1985;
    if(destProcID == 38) return 1986;
    if(destProcID == 45) return 1987;
    if(destProcID == 51) return 1988;
    if(destProcID == 61) return 1989;
    if(destProcID == 66) return 1990;
    if(destProcID == 89) return 1991;
    if(destProcID == 87) return 1992;
    if(destProcID == 78) return 1993;
    if(destProcID == 70) return 1994;
    if(destProcID == 56) return 1995;
    if(destProcID == 52) return 1996;
    if(destProcID == 9) return 1997;
    if(destProcID == 2) return 1998;
    if(destProcID == 129) return 1999;
    if(destProcID == 119) return 2000;
    if(destProcID == 114) return 2001;
  end
  if (srcProcId == 91) begin
    if(destProcID == 92) return 2002;
    if(destProcID == 94) return 2003;
    if(destProcID == 103) return 2004;
    if(destProcID == 111) return 2005;
    if(destProcID == 125) return 2006;
    if(destProcID == 129) return 2007;
    if(destProcID == 39) return 2008;
    if(destProcID == 46) return 2009;
    if(destProcID == 52) return 2010;
    if(destProcID == 62) return 2011;
    if(destProcID == 67) return 2012;
    if(destProcID == 90) return 2013;
    if(destProcID == 88) return 2014;
    if(destProcID == 79) return 2015;
    if(destProcID == 71) return 2016;
    if(destProcID == 57) return 2017;
    if(destProcID == 53) return 2018;
    if(destProcID == 10) return 2019;
    if(destProcID == 3) return 2020;
    if(destProcID == 130) return 2021;
    if(destProcID == 120) return 2022;
    if(destProcID == 115) return 2023;
  end
  if (srcProcId == 92) begin
    if(destProcID == 93) return 2024;
    if(destProcID == 95) return 2025;
    if(destProcID == 104) return 2026;
    if(destProcID == 112) return 2027;
    if(destProcID == 126) return 2028;
    if(destProcID == 130) return 2029;
    if(destProcID == 40) return 2030;
    if(destProcID == 47) return 2031;
    if(destProcID == 53) return 2032;
    if(destProcID == 63) return 2033;
    if(destProcID == 68) return 2034;
    if(destProcID == 91) return 2035;
    if(destProcID == 89) return 2036;
    if(destProcID == 80) return 2037;
    if(destProcID == 72) return 2038;
    if(destProcID == 58) return 2039;
    if(destProcID == 54) return 2040;
    if(destProcID == 11) return 2041;
    if(destProcID == 4) return 2042;
    if(destProcID == 131) return 2043;
    if(destProcID == 121) return 2044;
    if(destProcID == 116) return 2045;
  end
  if (srcProcId == 93) begin
    if(destProcID == 94) return 2046;
    if(destProcID == 96) return 2047;
    if(destProcID == 105) return 2048;
    if(destProcID == 113) return 2049;
    if(destProcID == 127) return 2050;
    if(destProcID == 131) return 2051;
    if(destProcID == 41) return 2052;
    if(destProcID == 48) return 2053;
    if(destProcID == 54) return 2054;
    if(destProcID == 64) return 2055;
    if(destProcID == 69) return 2056;
    if(destProcID == 92) return 2057;
    if(destProcID == 90) return 2058;
    if(destProcID == 81) return 2059;
    if(destProcID == 73) return 2060;
    if(destProcID == 59) return 2061;
    if(destProcID == 55) return 2062;
    if(destProcID == 12) return 2063;
    if(destProcID == 5) return 2064;
    if(destProcID == 132) return 2065;
    if(destProcID == 122) return 2066;
    if(destProcID == 117) return 2067;
  end
  if (srcProcId == 94) begin
    if(destProcID == 95) return 2068;
    if(destProcID == 97) return 2069;
    if(destProcID == 106) return 2070;
    if(destProcID == 114) return 2071;
    if(destProcID == 128) return 2072;
    if(destProcID == 132) return 2073;
    if(destProcID == 42) return 2074;
    if(destProcID == 49) return 2075;
    if(destProcID == 55) return 2076;
    if(destProcID == 65) return 2077;
    if(destProcID == 70) return 2078;
    if(destProcID == 93) return 2079;
    if(destProcID == 91) return 2080;
    if(destProcID == 82) return 2081;
    if(destProcID == 74) return 2082;
    if(destProcID == 60) return 2083;
    if(destProcID == 56) return 2084;
    if(destProcID == 13) return 2085;
    if(destProcID == 6) return 2086;
    if(destProcID == 0) return 2087;
    if(destProcID == 123) return 2088;
    if(destProcID == 118) return 2089;
  end
  if (srcProcId == 95) begin
    if(destProcID == 96) return 2090;
    if(destProcID == 98) return 2091;
    if(destProcID == 107) return 2092;
    if(destProcID == 115) return 2093;
    if(destProcID == 129) return 2094;
    if(destProcID == 0) return 2095;
    if(destProcID == 43) return 2096;
    if(destProcID == 50) return 2097;
    if(destProcID == 56) return 2098;
    if(destProcID == 66) return 2099;
    if(destProcID == 71) return 2100;
    if(destProcID == 94) return 2101;
    if(destProcID == 92) return 2102;
    if(destProcID == 83) return 2103;
    if(destProcID == 75) return 2104;
    if(destProcID == 61) return 2105;
    if(destProcID == 57) return 2106;
    if(destProcID == 14) return 2107;
    if(destProcID == 7) return 2108;
    if(destProcID == 1) return 2109;
    if(destProcID == 124) return 2110;
    if(destProcID == 119) return 2111;
  end
  if (srcProcId == 96) begin
    if(destProcID == 97) return 2112;
    if(destProcID == 99) return 2113;
    if(destProcID == 108) return 2114;
    if(destProcID == 116) return 2115;
    if(destProcID == 130) return 2116;
    if(destProcID == 1) return 2117;
    if(destProcID == 44) return 2118;
    if(destProcID == 51) return 2119;
    if(destProcID == 57) return 2120;
    if(destProcID == 67) return 2121;
    if(destProcID == 72) return 2122;
    if(destProcID == 95) return 2123;
    if(destProcID == 93) return 2124;
    if(destProcID == 84) return 2125;
    if(destProcID == 76) return 2126;
    if(destProcID == 62) return 2127;
    if(destProcID == 58) return 2128;
    if(destProcID == 15) return 2129;
    if(destProcID == 8) return 2130;
    if(destProcID == 2) return 2131;
    if(destProcID == 125) return 2132;
    if(destProcID == 120) return 2133;
  end
  if (srcProcId == 97) begin
    if(destProcID == 98) return 2134;
    if(destProcID == 100) return 2135;
    if(destProcID == 109) return 2136;
    if(destProcID == 117) return 2137;
    if(destProcID == 131) return 2138;
    if(destProcID == 2) return 2139;
    if(destProcID == 45) return 2140;
    if(destProcID == 52) return 2141;
    if(destProcID == 58) return 2142;
    if(destProcID == 68) return 2143;
    if(destProcID == 73) return 2144;
    if(destProcID == 96) return 2145;
    if(destProcID == 94) return 2146;
    if(destProcID == 85) return 2147;
    if(destProcID == 77) return 2148;
    if(destProcID == 63) return 2149;
    if(destProcID == 59) return 2150;
    if(destProcID == 16) return 2151;
    if(destProcID == 9) return 2152;
    if(destProcID == 3) return 2153;
    if(destProcID == 126) return 2154;
    if(destProcID == 121) return 2155;
  end
  if (srcProcId == 98) begin
    if(destProcID == 99) return 2156;
    if(destProcID == 101) return 2157;
    if(destProcID == 110) return 2158;
    if(destProcID == 118) return 2159;
    if(destProcID == 132) return 2160;
    if(destProcID == 3) return 2161;
    if(destProcID == 46) return 2162;
    if(destProcID == 53) return 2163;
    if(destProcID == 59) return 2164;
    if(destProcID == 69) return 2165;
    if(destProcID == 74) return 2166;
    if(destProcID == 97) return 2167;
    if(destProcID == 95) return 2168;
    if(destProcID == 86) return 2169;
    if(destProcID == 78) return 2170;
    if(destProcID == 64) return 2171;
    if(destProcID == 60) return 2172;
    if(destProcID == 17) return 2173;
    if(destProcID == 10) return 2174;
    if(destProcID == 4) return 2175;
    if(destProcID == 127) return 2176;
    if(destProcID == 122) return 2177;
  end
  if (srcProcId == 99) begin
    if(destProcID == 100) return 2178;
    if(destProcID == 102) return 2179;
    if(destProcID == 111) return 2180;
    if(destProcID == 119) return 2181;
    if(destProcID == 0) return 2182;
    if(destProcID == 4) return 2183;
    if(destProcID == 47) return 2184;
    if(destProcID == 54) return 2185;
    if(destProcID == 60) return 2186;
    if(destProcID == 70) return 2187;
    if(destProcID == 75) return 2188;
    if(destProcID == 98) return 2189;
    if(destProcID == 96) return 2190;
    if(destProcID == 87) return 2191;
    if(destProcID == 79) return 2192;
    if(destProcID == 65) return 2193;
    if(destProcID == 61) return 2194;
    if(destProcID == 18) return 2195;
    if(destProcID == 11) return 2196;
    if(destProcID == 5) return 2197;
    if(destProcID == 128) return 2198;
    if(destProcID == 123) return 2199;
  end
  if (srcProcId == 100) begin
    if(destProcID == 101) return 2200;
    if(destProcID == 103) return 2201;
    if(destProcID == 112) return 2202;
    if(destProcID == 120) return 2203;
    if(destProcID == 1) return 2204;
    if(destProcID == 5) return 2205;
    if(destProcID == 48) return 2206;
    if(destProcID == 55) return 2207;
    if(destProcID == 61) return 2208;
    if(destProcID == 71) return 2209;
    if(destProcID == 76) return 2210;
    if(destProcID == 99) return 2211;
    if(destProcID == 97) return 2212;
    if(destProcID == 88) return 2213;
    if(destProcID == 80) return 2214;
    if(destProcID == 66) return 2215;
    if(destProcID == 62) return 2216;
    if(destProcID == 19) return 2217;
    if(destProcID == 12) return 2218;
    if(destProcID == 6) return 2219;
    if(destProcID == 129) return 2220;
    if(destProcID == 124) return 2221;
  end
  if (srcProcId == 101) begin
    if(destProcID == 102) return 2222;
    if(destProcID == 104) return 2223;
    if(destProcID == 113) return 2224;
    if(destProcID == 121) return 2225;
    if(destProcID == 2) return 2226;
    if(destProcID == 6) return 2227;
    if(destProcID == 49) return 2228;
    if(destProcID == 56) return 2229;
    if(destProcID == 62) return 2230;
    if(destProcID == 72) return 2231;
    if(destProcID == 77) return 2232;
    if(destProcID == 100) return 2233;
    if(destProcID == 98) return 2234;
    if(destProcID == 89) return 2235;
    if(destProcID == 81) return 2236;
    if(destProcID == 67) return 2237;
    if(destProcID == 63) return 2238;
    if(destProcID == 20) return 2239;
    if(destProcID == 13) return 2240;
    if(destProcID == 7) return 2241;
    if(destProcID == 130) return 2242;
    if(destProcID == 125) return 2243;
  end
  if (srcProcId == 102) begin
    if(destProcID == 103) return 2244;
    if(destProcID == 105) return 2245;
    if(destProcID == 114) return 2246;
    if(destProcID == 122) return 2247;
    if(destProcID == 3) return 2248;
    if(destProcID == 7) return 2249;
    if(destProcID == 50) return 2250;
    if(destProcID == 57) return 2251;
    if(destProcID == 63) return 2252;
    if(destProcID == 73) return 2253;
    if(destProcID == 78) return 2254;
    if(destProcID == 101) return 2255;
    if(destProcID == 99) return 2256;
    if(destProcID == 90) return 2257;
    if(destProcID == 82) return 2258;
    if(destProcID == 68) return 2259;
    if(destProcID == 64) return 2260;
    if(destProcID == 21) return 2261;
    if(destProcID == 14) return 2262;
    if(destProcID == 8) return 2263;
    if(destProcID == 131) return 2264;
    if(destProcID == 126) return 2265;
  end
  if (srcProcId == 103) begin
    if(destProcID == 104) return 2266;
    if(destProcID == 106) return 2267;
    if(destProcID == 115) return 2268;
    if(destProcID == 123) return 2269;
    if(destProcID == 4) return 2270;
    if(destProcID == 8) return 2271;
    if(destProcID == 51) return 2272;
    if(destProcID == 58) return 2273;
    if(destProcID == 64) return 2274;
    if(destProcID == 74) return 2275;
    if(destProcID == 79) return 2276;
    if(destProcID == 102) return 2277;
    if(destProcID == 100) return 2278;
    if(destProcID == 91) return 2279;
    if(destProcID == 83) return 2280;
    if(destProcID == 69) return 2281;
    if(destProcID == 65) return 2282;
    if(destProcID == 22) return 2283;
    if(destProcID == 15) return 2284;
    if(destProcID == 9) return 2285;
    if(destProcID == 132) return 2286;
    if(destProcID == 127) return 2287;
  end
  if (srcProcId == 104) begin
    if(destProcID == 105) return 2288;
    if(destProcID == 107) return 2289;
    if(destProcID == 116) return 2290;
    if(destProcID == 124) return 2291;
    if(destProcID == 5) return 2292;
    if(destProcID == 9) return 2293;
    if(destProcID == 52) return 2294;
    if(destProcID == 59) return 2295;
    if(destProcID == 65) return 2296;
    if(destProcID == 75) return 2297;
    if(destProcID == 80) return 2298;
    if(destProcID == 103) return 2299;
    if(destProcID == 101) return 2300;
    if(destProcID == 92) return 2301;
    if(destProcID == 84) return 2302;
    if(destProcID == 70) return 2303;
    if(destProcID == 66) return 2304;
    if(destProcID == 23) return 2305;
    if(destProcID == 16) return 2306;
    if(destProcID == 10) return 2307;
    if(destProcID == 0) return 2308;
    if(destProcID == 128) return 2309;
  end
  if (srcProcId == 105) begin
    if(destProcID == 106) return 2310;
    if(destProcID == 108) return 2311;
    if(destProcID == 117) return 2312;
    if(destProcID == 125) return 2313;
    if(destProcID == 6) return 2314;
    if(destProcID == 10) return 2315;
    if(destProcID == 53) return 2316;
    if(destProcID == 60) return 2317;
    if(destProcID == 66) return 2318;
    if(destProcID == 76) return 2319;
    if(destProcID == 81) return 2320;
    if(destProcID == 104) return 2321;
    if(destProcID == 102) return 2322;
    if(destProcID == 93) return 2323;
    if(destProcID == 85) return 2324;
    if(destProcID == 71) return 2325;
    if(destProcID == 67) return 2326;
    if(destProcID == 24) return 2327;
    if(destProcID == 17) return 2328;
    if(destProcID == 11) return 2329;
    if(destProcID == 1) return 2330;
    if(destProcID == 129) return 2331;
  end
  if (srcProcId == 106) begin
    if(destProcID == 107) return 2332;
    if(destProcID == 109) return 2333;
    if(destProcID == 118) return 2334;
    if(destProcID == 126) return 2335;
    if(destProcID == 7) return 2336;
    if(destProcID == 11) return 2337;
    if(destProcID == 54) return 2338;
    if(destProcID == 61) return 2339;
    if(destProcID == 67) return 2340;
    if(destProcID == 77) return 2341;
    if(destProcID == 82) return 2342;
    if(destProcID == 105) return 2343;
    if(destProcID == 103) return 2344;
    if(destProcID == 94) return 2345;
    if(destProcID == 86) return 2346;
    if(destProcID == 72) return 2347;
    if(destProcID == 68) return 2348;
    if(destProcID == 25) return 2349;
    if(destProcID == 18) return 2350;
    if(destProcID == 12) return 2351;
    if(destProcID == 2) return 2352;
    if(destProcID == 130) return 2353;
  end
  if (srcProcId == 107) begin
    if(destProcID == 108) return 2354;
    if(destProcID == 110) return 2355;
    if(destProcID == 119) return 2356;
    if(destProcID == 127) return 2357;
    if(destProcID == 8) return 2358;
    if(destProcID == 12) return 2359;
    if(destProcID == 55) return 2360;
    if(destProcID == 62) return 2361;
    if(destProcID == 68) return 2362;
    if(destProcID == 78) return 2363;
    if(destProcID == 83) return 2364;
    if(destProcID == 106) return 2365;
    if(destProcID == 104) return 2366;
    if(destProcID == 95) return 2367;
    if(destProcID == 87) return 2368;
    if(destProcID == 73) return 2369;
    if(destProcID == 69) return 2370;
    if(destProcID == 26) return 2371;
    if(destProcID == 19) return 2372;
    if(destProcID == 13) return 2373;
    if(destProcID == 3) return 2374;
    if(destProcID == 131) return 2375;
  end
  if (srcProcId == 108) begin
    if(destProcID == 109) return 2376;
    if(destProcID == 111) return 2377;
    if(destProcID == 120) return 2378;
    if(destProcID == 128) return 2379;
    if(destProcID == 9) return 2380;
    if(destProcID == 13) return 2381;
    if(destProcID == 56) return 2382;
    if(destProcID == 63) return 2383;
    if(destProcID == 69) return 2384;
    if(destProcID == 79) return 2385;
    if(destProcID == 84) return 2386;
    if(destProcID == 107) return 2387;
    if(destProcID == 105) return 2388;
    if(destProcID == 96) return 2389;
    if(destProcID == 88) return 2390;
    if(destProcID == 74) return 2391;
    if(destProcID == 70) return 2392;
    if(destProcID == 27) return 2393;
    if(destProcID == 20) return 2394;
    if(destProcID == 14) return 2395;
    if(destProcID == 4) return 2396;
    if(destProcID == 132) return 2397;
  end
  if (srcProcId == 109) begin
    if(destProcID == 110) return 2398;
    if(destProcID == 112) return 2399;
    if(destProcID == 121) return 2400;
    if(destProcID == 129) return 2401;
    if(destProcID == 10) return 2402;
    if(destProcID == 14) return 2403;
    if(destProcID == 57) return 2404;
    if(destProcID == 64) return 2405;
    if(destProcID == 70) return 2406;
    if(destProcID == 80) return 2407;
    if(destProcID == 85) return 2408;
    if(destProcID == 108) return 2409;
    if(destProcID == 106) return 2410;
    if(destProcID == 97) return 2411;
    if(destProcID == 89) return 2412;
    if(destProcID == 75) return 2413;
    if(destProcID == 71) return 2414;
    if(destProcID == 28) return 2415;
    if(destProcID == 21) return 2416;
    if(destProcID == 15) return 2417;
    if(destProcID == 5) return 2418;
    if(destProcID == 0) return 2419;
  end
  if (srcProcId == 110) begin
    if(destProcID == 111) return 2420;
    if(destProcID == 113) return 2421;
    if(destProcID == 122) return 2422;
    if(destProcID == 130) return 2423;
    if(destProcID == 11) return 2424;
    if(destProcID == 15) return 2425;
    if(destProcID == 58) return 2426;
    if(destProcID == 65) return 2427;
    if(destProcID == 71) return 2428;
    if(destProcID == 81) return 2429;
    if(destProcID == 86) return 2430;
    if(destProcID == 109) return 2431;
    if(destProcID == 107) return 2432;
    if(destProcID == 98) return 2433;
    if(destProcID == 90) return 2434;
    if(destProcID == 76) return 2435;
    if(destProcID == 72) return 2436;
    if(destProcID == 29) return 2437;
    if(destProcID == 22) return 2438;
    if(destProcID == 16) return 2439;
    if(destProcID == 6) return 2440;
    if(destProcID == 1) return 2441;
  end
  if (srcProcId == 111) begin
    if(destProcID == 112) return 2442;
    if(destProcID == 114) return 2443;
    if(destProcID == 123) return 2444;
    if(destProcID == 131) return 2445;
    if(destProcID == 12) return 2446;
    if(destProcID == 16) return 2447;
    if(destProcID == 59) return 2448;
    if(destProcID == 66) return 2449;
    if(destProcID == 72) return 2450;
    if(destProcID == 82) return 2451;
    if(destProcID == 87) return 2452;
    if(destProcID == 110) return 2453;
    if(destProcID == 108) return 2454;
    if(destProcID == 99) return 2455;
    if(destProcID == 91) return 2456;
    if(destProcID == 77) return 2457;
    if(destProcID == 73) return 2458;
    if(destProcID == 30) return 2459;
    if(destProcID == 23) return 2460;
    if(destProcID == 17) return 2461;
    if(destProcID == 7) return 2462;
    if(destProcID == 2) return 2463;
  end
  if (srcProcId == 112) begin
    if(destProcID == 113) return 2464;
    if(destProcID == 115) return 2465;
    if(destProcID == 124) return 2466;
    if(destProcID == 132) return 2467;
    if(destProcID == 13) return 2468;
    if(destProcID == 17) return 2469;
    if(destProcID == 60) return 2470;
    if(destProcID == 67) return 2471;
    if(destProcID == 73) return 2472;
    if(destProcID == 83) return 2473;
    if(destProcID == 88) return 2474;
    if(destProcID == 111) return 2475;
    if(destProcID == 109) return 2476;
    if(destProcID == 100) return 2477;
    if(destProcID == 92) return 2478;
    if(destProcID == 78) return 2479;
    if(destProcID == 74) return 2480;
    if(destProcID == 31) return 2481;
    if(destProcID == 24) return 2482;
    if(destProcID == 18) return 2483;
    if(destProcID == 8) return 2484;
    if(destProcID == 3) return 2485;
  end
  if (srcProcId == 113) begin
    if(destProcID == 114) return 2486;
    if(destProcID == 116) return 2487;
    if(destProcID == 125) return 2488;
    if(destProcID == 0) return 2489;
    if(destProcID == 14) return 2490;
    if(destProcID == 18) return 2491;
    if(destProcID == 61) return 2492;
    if(destProcID == 68) return 2493;
    if(destProcID == 74) return 2494;
    if(destProcID == 84) return 2495;
    if(destProcID == 89) return 2496;
    if(destProcID == 112) return 2497;
    if(destProcID == 110) return 2498;
    if(destProcID == 101) return 2499;
    if(destProcID == 93) return 2500;
    if(destProcID == 79) return 2501;
    if(destProcID == 75) return 2502;
    if(destProcID == 32) return 2503;
    if(destProcID == 25) return 2504;
    if(destProcID == 19) return 2505;
    if(destProcID == 9) return 2506;
    if(destProcID == 4) return 2507;
  end
  if (srcProcId == 114) begin
    if(destProcID == 115) return 2508;
    if(destProcID == 117) return 2509;
    if(destProcID == 126) return 2510;
    if(destProcID == 1) return 2511;
    if(destProcID == 15) return 2512;
    if(destProcID == 19) return 2513;
    if(destProcID == 62) return 2514;
    if(destProcID == 69) return 2515;
    if(destProcID == 75) return 2516;
    if(destProcID == 85) return 2517;
    if(destProcID == 90) return 2518;
    if(destProcID == 113) return 2519;
    if(destProcID == 111) return 2520;
    if(destProcID == 102) return 2521;
    if(destProcID == 94) return 2522;
    if(destProcID == 80) return 2523;
    if(destProcID == 76) return 2524;
    if(destProcID == 33) return 2525;
    if(destProcID == 26) return 2526;
    if(destProcID == 20) return 2527;
    if(destProcID == 10) return 2528;
    if(destProcID == 5) return 2529;
  end
  if (srcProcId == 115) begin
    if(destProcID == 116) return 2530;
    if(destProcID == 118) return 2531;
    if(destProcID == 127) return 2532;
    if(destProcID == 2) return 2533;
    if(destProcID == 16) return 2534;
    if(destProcID == 20) return 2535;
    if(destProcID == 63) return 2536;
    if(destProcID == 70) return 2537;
    if(destProcID == 76) return 2538;
    if(destProcID == 86) return 2539;
    if(destProcID == 91) return 2540;
    if(destProcID == 114) return 2541;
    if(destProcID == 112) return 2542;
    if(destProcID == 103) return 2543;
    if(destProcID == 95) return 2544;
    if(destProcID == 81) return 2545;
    if(destProcID == 77) return 2546;
    if(destProcID == 34) return 2547;
    if(destProcID == 27) return 2548;
    if(destProcID == 21) return 2549;
    if(destProcID == 11) return 2550;
    if(destProcID == 6) return 2551;
  end
  if (srcProcId == 116) begin
    if(destProcID == 117) return 2552;
    if(destProcID == 119) return 2553;
    if(destProcID == 128) return 2554;
    if(destProcID == 3) return 2555;
    if(destProcID == 17) return 2556;
    if(destProcID == 21) return 2557;
    if(destProcID == 64) return 2558;
    if(destProcID == 71) return 2559;
    if(destProcID == 77) return 2560;
    if(destProcID == 87) return 2561;
    if(destProcID == 92) return 2562;
    if(destProcID == 115) return 2563;
    if(destProcID == 113) return 2564;
    if(destProcID == 104) return 2565;
    if(destProcID == 96) return 2566;
    if(destProcID == 82) return 2567;
    if(destProcID == 78) return 2568;
    if(destProcID == 35) return 2569;
    if(destProcID == 28) return 2570;
    if(destProcID == 22) return 2571;
    if(destProcID == 12) return 2572;
    if(destProcID == 7) return 2573;
  end
  if (srcProcId == 117) begin
    if(destProcID == 118) return 2574;
    if(destProcID == 120) return 2575;
    if(destProcID == 129) return 2576;
    if(destProcID == 4) return 2577;
    if(destProcID == 18) return 2578;
    if(destProcID == 22) return 2579;
    if(destProcID == 65) return 2580;
    if(destProcID == 72) return 2581;
    if(destProcID == 78) return 2582;
    if(destProcID == 88) return 2583;
    if(destProcID == 93) return 2584;
    if(destProcID == 116) return 2585;
    if(destProcID == 114) return 2586;
    if(destProcID == 105) return 2587;
    if(destProcID == 97) return 2588;
    if(destProcID == 83) return 2589;
    if(destProcID == 79) return 2590;
    if(destProcID == 36) return 2591;
    if(destProcID == 29) return 2592;
    if(destProcID == 23) return 2593;
    if(destProcID == 13) return 2594;
    if(destProcID == 8) return 2595;
  end
  if (srcProcId == 118) begin
    if(destProcID == 119) return 2596;
    if(destProcID == 121) return 2597;
    if(destProcID == 130) return 2598;
    if(destProcID == 5) return 2599;
    if(destProcID == 19) return 2600;
    if(destProcID == 23) return 2601;
    if(destProcID == 66) return 2602;
    if(destProcID == 73) return 2603;
    if(destProcID == 79) return 2604;
    if(destProcID == 89) return 2605;
    if(destProcID == 94) return 2606;
    if(destProcID == 117) return 2607;
    if(destProcID == 115) return 2608;
    if(destProcID == 106) return 2609;
    if(destProcID == 98) return 2610;
    if(destProcID == 84) return 2611;
    if(destProcID == 80) return 2612;
    if(destProcID == 37) return 2613;
    if(destProcID == 30) return 2614;
    if(destProcID == 24) return 2615;
    if(destProcID == 14) return 2616;
    if(destProcID == 9) return 2617;
  end
  if (srcProcId == 119) begin
    if(destProcID == 120) return 2618;
    if(destProcID == 122) return 2619;
    if(destProcID == 131) return 2620;
    if(destProcID == 6) return 2621;
    if(destProcID == 20) return 2622;
    if(destProcID == 24) return 2623;
    if(destProcID == 67) return 2624;
    if(destProcID == 74) return 2625;
    if(destProcID == 80) return 2626;
    if(destProcID == 90) return 2627;
    if(destProcID == 95) return 2628;
    if(destProcID == 118) return 2629;
    if(destProcID == 116) return 2630;
    if(destProcID == 107) return 2631;
    if(destProcID == 99) return 2632;
    if(destProcID == 85) return 2633;
    if(destProcID == 81) return 2634;
    if(destProcID == 38) return 2635;
    if(destProcID == 31) return 2636;
    if(destProcID == 25) return 2637;
    if(destProcID == 15) return 2638;
    if(destProcID == 10) return 2639;
  end
  if (srcProcId == 120) begin
    if(destProcID == 121) return 2640;
    if(destProcID == 123) return 2641;
    if(destProcID == 132) return 2642;
    if(destProcID == 7) return 2643;
    if(destProcID == 21) return 2644;
    if(destProcID == 25) return 2645;
    if(destProcID == 68) return 2646;
    if(destProcID == 75) return 2647;
    if(destProcID == 81) return 2648;
    if(destProcID == 91) return 2649;
    if(destProcID == 96) return 2650;
    if(destProcID == 119) return 2651;
    if(destProcID == 117) return 2652;
    if(destProcID == 108) return 2653;
    if(destProcID == 100) return 2654;
    if(destProcID == 86) return 2655;
    if(destProcID == 82) return 2656;
    if(destProcID == 39) return 2657;
    if(destProcID == 32) return 2658;
    if(destProcID == 26) return 2659;
    if(destProcID == 16) return 2660;
    if(destProcID == 11) return 2661;
  end
  if (srcProcId == 121) begin
    if(destProcID == 122) return 2662;
    if(destProcID == 124) return 2663;
    if(destProcID == 0) return 2664;
    if(destProcID == 8) return 2665;
    if(destProcID == 22) return 2666;
    if(destProcID == 26) return 2667;
    if(destProcID == 69) return 2668;
    if(destProcID == 76) return 2669;
    if(destProcID == 82) return 2670;
    if(destProcID == 92) return 2671;
    if(destProcID == 97) return 2672;
    if(destProcID == 120) return 2673;
    if(destProcID == 118) return 2674;
    if(destProcID == 109) return 2675;
    if(destProcID == 101) return 2676;
    if(destProcID == 87) return 2677;
    if(destProcID == 83) return 2678;
    if(destProcID == 40) return 2679;
    if(destProcID == 33) return 2680;
    if(destProcID == 27) return 2681;
    if(destProcID == 17) return 2682;
    if(destProcID == 12) return 2683;
  end
  if (srcProcId == 122) begin
    if(destProcID == 123) return 2684;
    if(destProcID == 125) return 2685;
    if(destProcID == 1) return 2686;
    if(destProcID == 9) return 2687;
    if(destProcID == 23) return 2688;
    if(destProcID == 27) return 2689;
    if(destProcID == 70) return 2690;
    if(destProcID == 77) return 2691;
    if(destProcID == 83) return 2692;
    if(destProcID == 93) return 2693;
    if(destProcID == 98) return 2694;
    if(destProcID == 121) return 2695;
    if(destProcID == 119) return 2696;
    if(destProcID == 110) return 2697;
    if(destProcID == 102) return 2698;
    if(destProcID == 88) return 2699;
    if(destProcID == 84) return 2700;
    if(destProcID == 41) return 2701;
    if(destProcID == 34) return 2702;
    if(destProcID == 28) return 2703;
    if(destProcID == 18) return 2704;
    if(destProcID == 13) return 2705;
  end
  if (srcProcId == 123) begin
    if(destProcID == 124) return 2706;
    if(destProcID == 126) return 2707;
    if(destProcID == 2) return 2708;
    if(destProcID == 10) return 2709;
    if(destProcID == 24) return 2710;
    if(destProcID == 28) return 2711;
    if(destProcID == 71) return 2712;
    if(destProcID == 78) return 2713;
    if(destProcID == 84) return 2714;
    if(destProcID == 94) return 2715;
    if(destProcID == 99) return 2716;
    if(destProcID == 122) return 2717;
    if(destProcID == 120) return 2718;
    if(destProcID == 111) return 2719;
    if(destProcID == 103) return 2720;
    if(destProcID == 89) return 2721;
    if(destProcID == 85) return 2722;
    if(destProcID == 42) return 2723;
    if(destProcID == 35) return 2724;
    if(destProcID == 29) return 2725;
    if(destProcID == 19) return 2726;
    if(destProcID == 14) return 2727;
  end
  if (srcProcId == 124) begin
    if(destProcID == 125) return 2728;
    if(destProcID == 127) return 2729;
    if(destProcID == 3) return 2730;
    if(destProcID == 11) return 2731;
    if(destProcID == 25) return 2732;
    if(destProcID == 29) return 2733;
    if(destProcID == 72) return 2734;
    if(destProcID == 79) return 2735;
    if(destProcID == 85) return 2736;
    if(destProcID == 95) return 2737;
    if(destProcID == 100) return 2738;
    if(destProcID == 123) return 2739;
    if(destProcID == 121) return 2740;
    if(destProcID == 112) return 2741;
    if(destProcID == 104) return 2742;
    if(destProcID == 90) return 2743;
    if(destProcID == 86) return 2744;
    if(destProcID == 43) return 2745;
    if(destProcID == 36) return 2746;
    if(destProcID == 30) return 2747;
    if(destProcID == 20) return 2748;
    if(destProcID == 15) return 2749;
  end
  if (srcProcId == 125) begin
    if(destProcID == 126) return 2750;
    if(destProcID == 128) return 2751;
    if(destProcID == 4) return 2752;
    if(destProcID == 12) return 2753;
    if(destProcID == 26) return 2754;
    if(destProcID == 30) return 2755;
    if(destProcID == 73) return 2756;
    if(destProcID == 80) return 2757;
    if(destProcID == 86) return 2758;
    if(destProcID == 96) return 2759;
    if(destProcID == 101) return 2760;
    if(destProcID == 124) return 2761;
    if(destProcID == 122) return 2762;
    if(destProcID == 113) return 2763;
    if(destProcID == 105) return 2764;
    if(destProcID == 91) return 2765;
    if(destProcID == 87) return 2766;
    if(destProcID == 44) return 2767;
    if(destProcID == 37) return 2768;
    if(destProcID == 31) return 2769;
    if(destProcID == 21) return 2770;
    if(destProcID == 16) return 2771;
  end
  if (srcProcId == 126) begin
    if(destProcID == 127) return 2772;
    if(destProcID == 129) return 2773;
    if(destProcID == 5) return 2774;
    if(destProcID == 13) return 2775;
    if(destProcID == 27) return 2776;
    if(destProcID == 31) return 2777;
    if(destProcID == 74) return 2778;
    if(destProcID == 81) return 2779;
    if(destProcID == 87) return 2780;
    if(destProcID == 97) return 2781;
    if(destProcID == 102) return 2782;
    if(destProcID == 125) return 2783;
    if(destProcID == 123) return 2784;
    if(destProcID == 114) return 2785;
    if(destProcID == 106) return 2786;
    if(destProcID == 92) return 2787;
    if(destProcID == 88) return 2788;
    if(destProcID == 45) return 2789;
    if(destProcID == 38) return 2790;
    if(destProcID == 32) return 2791;
    if(destProcID == 22) return 2792;
    if(destProcID == 17) return 2793;
  end
  if (srcProcId == 127) begin
    if(destProcID == 128) return 2794;
    if(destProcID == 130) return 2795;
    if(destProcID == 6) return 2796;
    if(destProcID == 14) return 2797;
    if(destProcID == 28) return 2798;
    if(destProcID == 32) return 2799;
    if(destProcID == 75) return 2800;
    if(destProcID == 82) return 2801;
    if(destProcID == 88) return 2802;
    if(destProcID == 98) return 2803;
    if(destProcID == 103) return 2804;
    if(destProcID == 126) return 2805;
    if(destProcID == 124) return 2806;
    if(destProcID == 115) return 2807;
    if(destProcID == 107) return 2808;
    if(destProcID == 93) return 2809;
    if(destProcID == 89) return 2810;
    if(destProcID == 46) return 2811;
    if(destProcID == 39) return 2812;
    if(destProcID == 33) return 2813;
    if(destProcID == 23) return 2814;
    if(destProcID == 18) return 2815;
  end
  if (srcProcId == 128) begin
    if(destProcID == 129) return 2816;
    if(destProcID == 131) return 2817;
    if(destProcID == 7) return 2818;
    if(destProcID == 15) return 2819;
    if(destProcID == 29) return 2820;
    if(destProcID == 33) return 2821;
    if(destProcID == 76) return 2822;
    if(destProcID == 83) return 2823;
    if(destProcID == 89) return 2824;
    if(destProcID == 99) return 2825;
    if(destProcID == 104) return 2826;
    if(destProcID == 127) return 2827;
    if(destProcID == 125) return 2828;
    if(destProcID == 116) return 2829;
    if(destProcID == 108) return 2830;
    if(destProcID == 94) return 2831;
    if(destProcID == 90) return 2832;
    if(destProcID == 47) return 2833;
    if(destProcID == 40) return 2834;
    if(destProcID == 34) return 2835;
    if(destProcID == 24) return 2836;
    if(destProcID == 19) return 2837;
  end
  if (srcProcId == 129) begin
    if(destProcID == 130) return 2838;
    if(destProcID == 132) return 2839;
    if(destProcID == 8) return 2840;
    if(destProcID == 16) return 2841;
    if(destProcID == 30) return 2842;
    if(destProcID == 34) return 2843;
    if(destProcID == 77) return 2844;
    if(destProcID == 84) return 2845;
    if(destProcID == 90) return 2846;
    if(destProcID == 100) return 2847;
    if(destProcID == 105) return 2848;
    if(destProcID == 128) return 2849;
    if(destProcID == 126) return 2850;
    if(destProcID == 117) return 2851;
    if(destProcID == 109) return 2852;
    if(destProcID == 95) return 2853;
    if(destProcID == 91) return 2854;
    if(destProcID == 48) return 2855;
    if(destProcID == 41) return 2856;
    if(destProcID == 35) return 2857;
    if(destProcID == 25) return 2858;
    if(destProcID == 20) return 2859;
  end
  if (srcProcId == 130) begin
    if(destProcID == 131) return 2860;
    if(destProcID == 0) return 2861;
    if(destProcID == 9) return 2862;
    if(destProcID == 17) return 2863;
    if(destProcID == 31) return 2864;
    if(destProcID == 35) return 2865;
    if(destProcID == 78) return 2866;
    if(destProcID == 85) return 2867;
    if(destProcID == 91) return 2868;
    if(destProcID == 101) return 2869;
    if(destProcID == 106) return 2870;
    if(destProcID == 129) return 2871;
    if(destProcID == 127) return 2872;
    if(destProcID == 118) return 2873;
    if(destProcID == 110) return 2874;
    if(destProcID == 96) return 2875;
    if(destProcID == 92) return 2876;
    if(destProcID == 49) return 2877;
    if(destProcID == 42) return 2878;
    if(destProcID == 36) return 2879;
    if(destProcID == 26) return 2880;
    if(destProcID == 21) return 2881;
  end
  if (srcProcId == 131) begin
    if(destProcID == 132) return 2882;
    if(destProcID == 1) return 2883;
    if(destProcID == 10) return 2884;
    if(destProcID == 18) return 2885;
    if(destProcID == 32) return 2886;
    if(destProcID == 36) return 2887;
    if(destProcID == 79) return 2888;
    if(destProcID == 86) return 2889;
    if(destProcID == 92) return 2890;
    if(destProcID == 102) return 2891;
    if(destProcID == 107) return 2892;
    if(destProcID == 130) return 2893;
    if(destProcID == 128) return 2894;
    if(destProcID == 119) return 2895;
    if(destProcID == 111) return 2896;
    if(destProcID == 97) return 2897;
    if(destProcID == 93) return 2898;
    if(destProcID == 50) return 2899;
    if(destProcID == 43) return 2900;
    if(destProcID == 37) return 2901;
    if(destProcID == 27) return 2902;
    if(destProcID == 22) return 2903;
  end
  if (srcProcId == 132) begin
    if(destProcID == 0) return 2904;
    if(destProcID == 2) return 2905;
    if(destProcID == 11) return 2906;
    if(destProcID == 19) return 2907;
    if(destProcID == 33) return 2908;
    if(destProcID == 37) return 2909;
    if(destProcID == 80) return 2910;
    if(destProcID == 87) return 2911;
    if(destProcID == 93) return 2912;
    if(destProcID == 103) return 2913;
    if(destProcID == 108) return 2914;
    if(destProcID == 131) return 2915;
    if(destProcID == 129) return 2916;
    if(destProcID == 120) return 2917;
    if(destProcID == 112) return 2918;
    if(destProcID == 98) return 2919;
    if(destProcID == 94) return 2920;
    if(destProcID == 51) return 2921;
    if(destProcID == 44) return 2922;
    if(destProcID == 38) return 2923;
    if(destProcID == 28) return 2924;
    if(destProcID == 23) return 2925;
  end
  if (srcProcId == 133) begin
  end
  if (srcProcId == 134) begin
  end
  if (srcProcId == 135) begin
  end
  if (srcProcId == 136) begin
  end
  if (srcProcId == 137) begin
  end
  if (srcProcId == 138) begin
  end
  if (srcProcId == 139) begin
  end
  if (srcProcId == 140) begin
  end
  if (srcProcId == 141) begin
  end
  if (srcProcId == 142) begin
  end
  if (srcProcId == 143) begin
  end
  else return 0;
endfunction


// Lookup function for destination node at each mesh node corresponding to the arc id and source mesh 
function String lookupArcDest ( NoCAddr2D thisRowAddr, NoCAddr2D thisColAddr, NoCArcId arc_index); 
endfunction 
  if ((thisRowAddr == 5) & (thisColAddr == 6)) begin 
    if (arc_index == 0) return "W"  ;
    if (arc_index == 1) return "W"  ;
    if (arc_index == 2) return "E"  ;
    if (arc_index == 3) return "E"  ;
    if (arc_index == 4) return "E"  ;
    if (arc_index == 5) return "E"  ;
    if (arc_index == 6) return "E"  ;
    if (arc_index == 7) return "W"  ;
    if (arc_index == 8) return "E"  ;
    if (arc_index == 9) return "E"  ;
    if (arc_index == 10) return "E"  ;
    if (arc_index == 11) return "E"  ;
    if (arc_index == 12) return "E"  ;
    if (arc_index == 13) return "W"  ;
    if (arc_index == 14) return "W"  ;
    if (arc_index == 15) return "E"  ;
    if (arc_index == 16) return "E"  ;
    if (arc_index == 17) return "E"  ;
    if (arc_index == 18) return "W"  ;
    if (arc_index == 19) return "W"  ;
    if (arc_index == 20) return "W"  ;
    if (arc_index == 21) return "E"  ;
    if (arc_index == 30) return "E"  ;
    if (arc_index == 33) return "H"  ;
    if (arc_index == 78) return "H"  ;
    if (arc_index == 84) return "E"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 113) return "E"  ;
    if (arc_index == 125) return "E"  ;
    if (arc_index == 128) return "E"  ;
    if (arc_index == 158) return "W"  ;
    if (arc_index == 159) return "W"  ;
    if (arc_index == 160) return "W"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 170) return "W"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 210) return "W"  ;
    if (arc_index == 212) return "W"  ;
    if (arc_index == 233) return "W"  ;
    if (arc_index == 265) return "W"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 269) return "W"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 277) return "H"  ;
    if (arc_index == 285) return "H"  ;
    if (arc_index == 296) return "W"  ;
    if (arc_index == 308) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 315) return "W"  ;
    if (arc_index == 327) return "W"  ;
    if (arc_index == 332) return "E"  ;
    if (arc_index == 340) return "E"  ;
    if (arc_index == 344) return "E"  ;
    if (arc_index == 356) return "E"  ;
    if (arc_index == 399) return "E"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 426) return "E"  ;
    if (arc_index == 436) return "E"  ;
    if (arc_index == 454) return "H"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 535) return "W"  ;
    if (arc_index == 538) return "H"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 603) return "W"  ;
    if (arc_index == 609) return "W"  ;
    if (arc_index == 610) return "W"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 642) return "W"  ;
    if (arc_index == 647) return "H"  ;
    if (arc_index == 649) return "H"  ;
    if (arc_index == 653) return "E"  ;
    if (arc_index == 654) return "W"  ;
    if (arc_index == 655) return "W"  ;
    if (arc_index == 663) return "W"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 686) return "W"  ;
    if (arc_index == 691) return "W"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 763) return "H"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 784) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 836) return "E"  ;
    if (arc_index == 839) return "E"  ;
    if (arc_index == 850) return "E"  ;
    if (arc_index == 851) return "E"  ;
    if (arc_index == 852) return "H"  ;
    if (arc_index == 863) return "H"  ;
    if (arc_index == 866) return "H"  ;
    if (arc_index == 869) return "H"  ;
    if (arc_index == 898) return "H"  ;
    if (arc_index == 905) return "H"  ;
    if (arc_index == 917) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 971) return "E"  ;
    if (arc_index == 991) return "E"  ;
    if (arc_index == 997) return "H"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1035) return "E"  ;
    if (arc_index == 1038) return "E"  ;
    if (arc_index == 1056) return "E"  ;
    if (arc_index == 1061) return "W"  ;
    if (arc_index == 1062) return "W"  ;
    if (arc_index == 1063) return "W"  ;
    if (arc_index == 1068) return "W"  ;
    if (arc_index == 1075) return "W"  ;
    if (arc_index == 1077) return "W"  ;
    if (arc_index == 1085) return "W"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1089) return "E"  ;
    if (arc_index == 1093) return "E"  ;
    if (arc_index == 1100) return "E"  ;
    if (arc_index == 1101) return "E"  ;
    if (arc_index == 1102) return "E"  ;
    if (arc_index == 1107) return "E"  ;
    if (arc_index == 1109) return "E"  ;
    if (arc_index == 1112) return "E"  ;
    if (arc_index == 1114) return "E"  ;
    if (arc_index == 1115) return "E"  ;
    if (arc_index == 1116) return "E"  ;
    if (arc_index == 1117) return "E"  ;
    if (arc_index == 1119) return "E"  ;
    if (arc_index == 1124) return "E"  ;
    if (arc_index == 1133) return "E"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1148) return "W"  ;
    if (arc_index == 1150) return "H"  ;
    if (arc_index == 1170) return "W"  ;
    if (arc_index == 1174) return "W"  ;
    if (arc_index == 1178) return "W"  ;
    if (arc_index == 1187) return "W"  ;
    if (arc_index == 1195) return "W"  ;
    if (arc_index == 1212) return "W"  ;
    if (arc_index == 1220) return "W"  ;
    if (arc_index == 1274) return "W"  ;
    if (arc_index == 1275) return "W"  ;
    if (arc_index == 1280) return "W"  ;
    if (arc_index == 1290) return "W"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1327) return "W"  ;
    if (arc_index == 1328) return "W"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1377) return "W"  ;
    if (arc_index == 1396) return "W"  ;
    if (arc_index == 1397) return "W"  ;
    if (arc_index == 1401) return "W"  ;
    if (arc_index == 1405) return "W"  ;
    if (arc_index == 1413) return "W"  ;
    if (arc_index == 1415) return "W"  ;
    if (arc_index == 1422) return "W"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1449) return "W"  ;
    if (arc_index == 1456) return "W"  ;
    if (arc_index == 1462) return "W"  ;
    if (arc_index == 1470) return "W"  ;
    if (arc_index == 1471) return "W"  ;
    if (arc_index == 1480) return "W"  ;
    if (arc_index == 1494) return "W"  ;
    if (arc_index == 1507) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1580) return "E"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1594) return "E"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1620) return "E"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1641) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1650) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1672) return "W"  ;
    if (arc_index == 1673) return "W"  ;
    if (arc_index == 1684) return "W"  ;
    if (arc_index == 1691) return "W"  ;
    if (arc_index == 1696) return "E"  ;
    if (arc_index == 1703) return "E"  ;
    if (arc_index == 1704) return "E"  ;
    if (arc_index == 1730) return "E"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1737) return "E"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1785) return "W"  ;
    if (arc_index == 1788) return "W"  ;
    if (arc_index == 1799) return "H"  ;
    if (arc_index == 1807) return "H"  ;
    if (arc_index == 1823) return "W"  ;
    if (arc_index == 1829) return "E"  ;
    if (arc_index == 1848) return "E"  ;
    if (arc_index == 1893) return "E"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 1901) return "E"  ;
    if (arc_index == 1903) return "E"  ;
    if (arc_index == 1907) return "E"  ;
    if (arc_index == 1908) return "E"  ;
    if (arc_index == 1922) return "E"  ;
    if (arc_index == 1936) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1953) return "E"  ;
    if (arc_index == 1954) return "H"  ;
    if (arc_index == 1966) return "H"  ;
    if (arc_index == 1979) return "H"  ;
    if (arc_index == 1982) return "H"  ;
    if (arc_index == 1988) return "H"  ;
    if (arc_index == 1994) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2036) return "E"  ;
    if (arc_index == 2042) return "E"  ;
    if (arc_index == 2053) return "E"  ;
    if (arc_index == 2087) return "H"  ;
    if (arc_index == 2090) return "W"  ;
    if (arc_index == 2095) return "H"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2182) return "H"  ;
    if (arc_index == 2220) return "H"  ;
    if (arc_index == 2237) return "H"  ;
    if (arc_index == 2247) return "W"  ;
    if (arc_index == 2249) return "E"  ;
    if (arc_index == 2250) return "E"  ;
    if (arc_index == 2252) return "E"  ;
    if (arc_index == 2253) return "W"  ;
    if (arc_index == 2254) return "W"  ;
    if (arc_index == 2257) return "W"  ;
    if (arc_index == 2258) return "E"  ;
    if (arc_index == 2260) return "E"  ;
    if (arc_index == 2262) return "E"  ;
    if (arc_index == 2264) return "W"  ;
    if (arc_index == 2265) return "W"  ;
    if (arc_index == 2274) return "W"  ;
    if (arc_index == 2280) return "W"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2308) return "H"  ;
    if (arc_index == 2320) return "H"  ;
    if (arc_index == 2331) return "H"  ;
    if (arc_index == 2346) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2419) return "H"  ;
    if (arc_index == 2449) return "H"  ;
    if (arc_index == 2451) return "E"  ;
    if (arc_index == 2489) return "H"  ;
    if (arc_index == 2507) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2537) return "E"  ;
    if (arc_index == 2543) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2614) return "E"  ;
    if (arc_index == 2620) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2664) return "H"  ;
    if (arc_index == 2670) return "E"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2689) return "E"  ;
    if (arc_index == 2690) return "E"  ;
    if (arc_index == 2696) return "E"  ;
    if (arc_index == 2705) return "E"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2738) return "W"  ;
    if (arc_index == 2749) return "W"  ;
    if (arc_index == 2782) return "W"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2861) return "H"  ;
    if (arc_index == 2867) return "H"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2894) return "E"  ;
    if (arc_index == 2895) return "E"  ;
    if (arc_index == 2902) return "E"  ;
    if (arc_index == 2904) return "H"  ;
    if (arc_index == 2912) return "W"  ;
    if (arc_index == 2915) return "W"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 4)) begin 
    if (arc_index == 0) return "H"  ;
    if (arc_index == 22) return "H"  ;
    if (arc_index == 23) return "E"  ;
    if (arc_index == 24) return "E"  ;
    if (arc_index == 25) return "E"  ;
    if (arc_index == 26) return "E"  ;
    if (arc_index == 27) return "E"  ;
    if (arc_index == 28) return "E"  ;
    if (arc_index == 29) return "E"  ;
    if (arc_index == 30) return "E"  ;
    if (arc_index == 31) return "E"  ;
    if (arc_index == 32) return "W"  ;
    if (arc_index == 33) return "E"  ;
    if (arc_index == 34) return "E"  ;
    if (arc_index == 35) return "E"  ;
    if (arc_index == 36) return "E"  ;
    if (arc_index == 37) return "E"  ;
    if (arc_index == 38) return "E"  ;
    if (arc_index == 39) return "E"  ;
    if (arc_index == 40) return "E"  ;
    if (arc_index == 41) return "E"  ;
    if (arc_index == 42) return "W"  ;
    if (arc_index == 43) return "E"  ;
    if (arc_index == 45) return "E"  ;
    if (arc_index == 48) return "E"  ;
    if (arc_index == 54) return "E"  ;
    if (arc_index == 55) return "H"  ;
    if (arc_index == 60) return "H"  ;
    if (arc_index == 66) return "H"  ;
    if (arc_index == 74) return "H"  ;
    if (arc_index == 96) return "H"  ;
    if (arc_index == 100) return "H"  ;
    if (arc_index == 117) return "H"  ;
    if (arc_index == 122) return "H"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 136) return "E"  ;
    if (arc_index == 138) return "E"  ;
    if (arc_index == 142) return "E"  ;
    if (arc_index == 148) return "E"  ;
    if (arc_index == 152) return "E"  ;
    if (arc_index == 180) return "E"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 210) return "W"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 229) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 279) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 299) return "H"  ;
    if (arc_index == 346) return "W"  ;
    if (arc_index == 371) return "W"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 404) return "W"  ;
    if (arc_index == 410) return "W"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 445) return "E"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 461) return "E"  ;
    if (arc_index == 476) return "H"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 560) return "H"  ;
    if (arc_index == 640) return "W"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 663) return "W"  ;
    if (arc_index == 669) return "H"  ;
    if (arc_index == 752) return "H"  ;
    if (arc_index == 779) return "H"  ;
    if (arc_index == 785) return "H"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 807) return "E"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 874) return "H"  ;
    if (arc_index == 888) return "H"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 895) return "E"  ;
    if (arc_index == 903) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 946) return "E"  ;
    if (arc_index == 978) return "W"  ;
    if (arc_index == 979) return "W"  ;
    if (arc_index == 993) return "E"  ;
    if (arc_index == 996) return "E"  ;
    if (arc_index == 997) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1008) return "E"  ;
    if (arc_index == 1009) return "E"  ;
    if (arc_index == 1014) return "E"  ;
    if (arc_index == 1019) return "H"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1041) return "E"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1166) return "W"  ;
    if (arc_index == 1169) return "W"  ;
    if (arc_index == 1172) return "H"  ;
    if (arc_index == 1179) return "W"  ;
    if (arc_index == 1184) return "W"  ;
    if (arc_index == 1189) return "E"  ;
    if (arc_index == 1194) return "E"  ;
    if (arc_index == 1199) return "E"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1207) return "E"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1211) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1214) return "E"  ;
    if (arc_index == 1215) return "E"  ;
    if (arc_index == 1217) return "E"  ;
    if (arc_index == 1218) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1230) return "E"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1266) return "W"  ;
    if (arc_index == 1288) return "W"  ;
    if (arc_index == 1293) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1390) return "W"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1439) return "W"  ;
    if (arc_index == 1448) return "W"  ;
    if (arc_index == 1462) return "W"  ;
    if (arc_index == 1470) return "W"  ;
    if (arc_index == 1499) return "W"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1522) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1611) return "E"  ;
    if (arc_index == 1627) return "E"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1697) return "E"  ;
    if (arc_index == 1698) return "E"  ;
    if (arc_index == 1723) return "E"  ;
    if (arc_index == 1731) return "E"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1775) return "E"  ;
    if (arc_index == 1776) return "E"  ;
    if (arc_index == 1802) return "W"  ;
    if (arc_index == 1821) return "H"  ;
    if (arc_index == 1834) return "E"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1856) return "E"  ;
    if (arc_index == 1864) return "W"  ;
    if (arc_index == 1923) return "E"  ;
    if (arc_index == 1929) return "E"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 1973) return "W"  ;
    if (arc_index == 1976) return "H"  ;
    if (arc_index == 1980) return "H"  ;
    if (arc_index == 1983) return "W"  ;
    if (arc_index == 2004) return "E"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2056) return "W"  ;
    if (arc_index == 2062) return "W"  ;
    if (arc_index == 2064) return "E"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2109) return "H"  ;
    if (arc_index == 2117) return "H"  ;
    if (arc_index == 2138) return "H"  ;
    if (arc_index == 2139) return "H"  ;
    if (arc_index == 2141) return "E"  ;
    if (arc_index == 2144) return "E"  ;
    if (arc_index == 2145) return "E"  ;
    if (arc_index == 2148) return "E"  ;
    if (arc_index == 2149) return "E"  ;
    if (arc_index == 2152) return "E"  ;
    if (arc_index == 2153) return "E"  ;
    if (arc_index == 2154) return "E"  ;
    if (arc_index == 2155) return "E"  ;
    if (arc_index == 2163) return "E"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2167) return "E"  ;
    if (arc_index == 2175) return "E"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2204) return "H"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2279) return "E"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2330) return "H"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2398) return "W"  ;
    if (arc_index == 2420) return "W"  ;
    if (arc_index == 2425) return "W"  ;
    if (arc_index == 2426) return "E"  ;
    if (arc_index == 2427) return "E"  ;
    if (arc_index == 2428) return "E"  ;
    if (arc_index == 2430) return "E"  ;
    if (arc_index == 2431) return "E"  ;
    if (arc_index == 2435) return "E"  ;
    if (arc_index == 2437) return "E"  ;
    if (arc_index == 2439) return "E"  ;
    if (arc_index == 2441) return "H"  ;
    if (arc_index == 2445) return "H"  ;
    if (arc_index == 2451) return "H"  ;
    if (arc_index == 2452) return "W"  ;
    if (arc_index == 2457) return "W"  ;
    if (arc_index == 2458) return "W"  ;
    if (arc_index == 2460) return "W"  ;
    if (arc_index == 2463) return "W"  ;
    if (arc_index == 2475) return "W"  ;
    if (arc_index == 2498) return "W"  ;
    if (arc_index == 2510) return "W"  ;
    if (arc_index == 2511) return "H"  ;
    if (arc_index == 2518) return "H"  ;
    if (arc_index == 2519) return "H"  ;
    if (arc_index == 2521) return "E"  ;
    if (arc_index == 2524) return "E"  ;
    if (arc_index == 2541) return "W"  ;
    if (arc_index == 2551) return "W"  ;
    if (arc_index == 2584) return "W"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2672) return "E"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2686) return "H"  ;
    if (arc_index == 2704) return "E"  ;
    if (arc_index == 2733) return "E"  ;
    if (arc_index == 2774) return "E"  ;
    if (arc_index == 2781) return "E"  ;
    if (arc_index == 2785) return "W"  ;
    if (arc_index == 2812) return "W"  ;
    if (arc_index == 2883) return "H"  ;
    if (arc_index == 2885) return "H"  ;
    if (arc_index == 2896) return "H"  ;
    if (arc_index == 2897) return "H"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 4)) begin 
    if (arc_index == 1) return "W"  ;
    if (arc_index == 3) return "W"  ;
    if (arc_index == 22) return "H"  ;
    if (arc_index == 25) return "H"  ;
    if (arc_index == 26) return "H"  ;
    if (arc_index == 28) return "H"  ;
    if (arc_index == 34) return "H"  ;
    if (arc_index == 35) return "W"  ;
    if (arc_index == 38) return "E"  ;
    if (arc_index == 41) return "W"  ;
    if (arc_index == 44) return "W"  ;
    if (arc_index == 45) return "W"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 47) return "W"  ;
    if (arc_index == 48) return "W"  ;
    if (arc_index == 49) return "W"  ;
    if (arc_index == 50) return "W"  ;
    if (arc_index == 51) return "W"  ;
    if (arc_index == 52) return "E"  ;
    if (arc_index == 53) return "E"  ;
    if (arc_index == 54) return "E"  ;
    if (arc_index == 55) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 57) return "E"  ;
    if (arc_index == 58) return "E"  ;
    if (arc_index == 59) return "W"  ;
    if (arc_index == 60) return "W"  ;
    if (arc_index == 61) return "W"  ;
    if (arc_index == 62) return "E"  ;
    if (arc_index == 63) return "E"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 65) return "E"  ;
    if (arc_index == 68) return "E"  ;
    if (arc_index == 72) return "E"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 77) return "H"  ;
    if (arc_index == 87) return "H"  ;
    if (arc_index == 96) return "W"  ;
    if (arc_index == 106) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 117) return "W"  ;
    if (arc_index == 122) return "H"  ;
    if (arc_index == 136) return "H"  ;
    if (arc_index == 138) return "W"  ;
    if (arc_index == 142) return "W"  ;
    if (arc_index == 148) return "W"  ;
    if (arc_index == 152) return "W"  ;
    if (arc_index == 159) return "W"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 222) return "W"  ;
    if (arc_index == 227) return "W"  ;
    if (arc_index == 238) return "W"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 321) return "H"  ;
    if (arc_index == 343) return "W"  ;
    if (arc_index == 346) return "W"  ;
    if (arc_index == 349) return "W"  ;
    if (arc_index == 362) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 386) return "W"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 410) return "W"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 445) return "W"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 458) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 474) return "E"  ;
    if (arc_index == 476) return "E"  ;
    if (arc_index == 490) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 497) return "E"  ;
    if (arc_index == 498) return "H"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 530) return "W"  ;
    if (arc_index == 540) return "W"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 582) return "H"  ;
    if (arc_index == 591) return "E"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 663) return "E"  ;
    if (arc_index == 674) return "E"  ;
    if (arc_index == 691) return "H"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 752) return "W"  ;
    if (arc_index == 785) return "W"  ;
    if (arc_index == 807) return "H"  ;
    if (arc_index == 812) return "E"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 888) return "W"  ;
    if (arc_index == 891) return "W"  ;
    if (arc_index == 895) return "W"  ;
    if (arc_index == 896) return "H"  ;
    if (arc_index == 903) return "H"  ;
    if (arc_index == 910) return "H"  ;
    if (arc_index == 923) return "E"  ;
    if (arc_index == 928) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 946) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 972) return "E"  ;
    if (arc_index == 987) return "E"  ;
    if (arc_index == 996) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1008) return "E"  ;
    if (arc_index == 1009) return "E"  ;
    if (arc_index == 1041) return "H"  ;
    if (arc_index == 1047) return "H"  ;
    if (arc_index == 1169) return "H"  ;
    if (arc_index == 1194) return "H"  ;
    if (arc_index == 1195) return "E"  ;
    if (arc_index == 1196) return "E"  ;
    if (arc_index == 1207) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1214) return "E"  ;
    if (arc_index == 1215) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1230) return "E"  ;
    if (arc_index == 1292) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1325) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1390) return "W"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1437) return "W"  ;
    if (arc_index == 1438) return "W"  ;
    if (arc_index == 1440) return "W"  ;
    if (arc_index == 1444) return "W"  ;
    if (arc_index == 1448) return "W"  ;
    if (arc_index == 1462) return "W"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1499) return "W"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1564) return "E"  ;
    if (arc_index == 1611) return "E"  ;
    if (arc_index == 1627) return "E"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1648) return "E"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1697) return "E"  ;
    if (arc_index == 1698) return "E"  ;
    if (arc_index == 1731) return "E"  ;
    if (arc_index == 1775) return "E"  ;
    if (arc_index == 1776) return "E"  ;
    if (arc_index == 1802) return "E"  ;
    if (arc_index == 1834) return "E"  ;
    if (arc_index == 1843) return "H"  ;
    if (arc_index == 1856) return "H"  ;
    if (arc_index == 1857) return "W"  ;
    if (arc_index == 1864) return "W"  ;
    if (arc_index == 1865) return "W"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1894) return "W"  ;
    if (arc_index == 1923) return "W"  ;
    if (arc_index == 1929) return "W"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 1972) return "W"  ;
    if (arc_index == 1980) return "W"  ;
    if (arc_index == 1983) return "W"  ;
    if (arc_index == 1998) return "H"  ;
    if (arc_index == 2006) return "H"  ;
    if (arc_index == 2012) return "H"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2048) return "E"  ;
    if (arc_index == 2054) return "W"  ;
    if (arc_index == 2056) return "W"  ;
    if (arc_index == 2061) return "E"  ;
    if (arc_index == 2062) return "E"  ;
    if (arc_index == 2064) return "E"  ;
    if (arc_index == 2067) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2091) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2131) return "H"  ;
    if (arc_index == 2138) return "H"  ;
    if (arc_index == 2139) return "H"  ;
    if (arc_index == 2144) return "H"  ;
    if (arc_index == 2145) return "E"  ;
    if (arc_index == 2148) return "E"  ;
    if (arc_index == 2149) return "E"  ;
    if (arc_index == 2152) return "E"  ;
    if (arc_index == 2153) return "W"  ;
    if (arc_index == 2154) return "W"  ;
    if (arc_index == 2155) return "W"  ;
    if (arc_index == 2156) return "E"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2163) return "E"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2167) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2169) return "E"  ;
    if (arc_index == 2174) return "E"  ;
    if (arc_index == 2175) return "E"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2189) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2226) return "H"  ;
    if (arc_index == 2275) return "W"  ;
    if (arc_index == 2281) return "W"  ;
    if (arc_index == 2283) return "W"  ;
    if (arc_index == 2352) return "H"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2424) return "W"  ;
    if (arc_index == 2425) return "E"  ;
    if (arc_index == 2445) return "E"  ;
    if (arc_index == 2451) return "E"  ;
    if (arc_index == 2457) return "E"  ;
    if (arc_index == 2458) return "E"  ;
    if (arc_index == 2463) return "H"  ;
    if (arc_index == 2475) return "H"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2510) return "E"  ;
    if (arc_index == 2518) return "E"  ;
    if (arc_index == 2519) return "E"  ;
    if (arc_index == 2533) return "H"  ;
    if (arc_index == 2541) return "H"  ;
    if (arc_index == 2551) return "H"  ;
    if (arc_index == 2580) return "E"  ;
    if (arc_index == 2584) return "E"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2665) return "W"  ;
    if (arc_index == 2680) return "W"  ;
    if (arc_index == 2686) return "W"  ;
    if (arc_index == 2704) return "W"  ;
    if (arc_index == 2708) return "H"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2774) return "W"  ;
    if (arc_index == 2781) return "W"  ;
    if (arc_index == 2785) return "W"  ;
    if (arc_index == 2789) return "W"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2883) return "E"  ;
    if (arc_index == 2885) return "E"  ;
    if (arc_index == 2896) return "E"  ;
    if (arc_index == 2897) return "E"  ;
    if (arc_index == 2905) return "H"  ;
    if (arc_index == 2919) return "W"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 2)) begin 
    if (arc_index == 1) return "H"  ;
    if (arc_index == 3) return "W"  ;
    if (arc_index == 44) return "H"  ;
    if (arc_index == 47) return "W"  ;
    if (arc_index == 59) return "W"  ;
    if (arc_index == 61) return "W"  ;
    if (arc_index == 66) return "E"  ;
    if (arc_index == 67) return "E"  ;
    if (arc_index == 68) return "E"  ;
    if (arc_index == 69) return "W"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 71) return "E"  ;
    if (arc_index == 72) return "E"  ;
    if (arc_index == 73) return "E"  ;
    if (arc_index == 74) return "E"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 76) return "E"  ;
    if (arc_index == 77) return "E"  ;
    if (arc_index == 78) return "E"  ;
    if (arc_index == 79) return "E"  ;
    if (arc_index == 80) return "E"  ;
    if (arc_index == 81) return "E"  ;
    if (arc_index == 82) return "E"  ;
    if (arc_index == 83) return "W"  ;
    if (arc_index == 84) return "E"  ;
    if (arc_index == 85) return "E"  ;
    if (arc_index == 86) return "E"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 99) return "H"  ;
    if (arc_index == 106) return "H"  ;
    if (arc_index == 107) return "H"  ;
    if (arc_index == 115) return "H"  ;
    if (arc_index == 138) return "H"  ;
    if (arc_index == 144) return "H"  ;
    if (arc_index == 145) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 222) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 343) return "H"  ;
    if (arc_index == 349) return "H"  ;
    if (arc_index == 380) return "E"  ;
    if (arc_index == 390) return "E"  ;
    if (arc_index == 395) return "E"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 442) return "W"  ;
    if (arc_index == 443) return "W"  ;
    if (arc_index == 444) return "W"  ;
    if (arc_index == 445) return "E"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 448) return "E"  ;
    if (arc_index == 454) return "E"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 456) return "E"  ;
    if (arc_index == 458) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 461) return "E"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 490) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 497) return "E"  ;
    if (arc_index == 498) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 520) return "H"  ;
    if (arc_index == 527) return "H"  ;
    if (arc_index == 530) return "H"  ;
    if (arc_index == 546) return "H"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 579) return "E"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 582) return "E"  ;
    if (arc_index == 591) return "E"  ;
    if (arc_index == 604) return "H"  ;
    if (arc_index == 640) return "H"  ;
    if (arc_index == 641) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 713) return "H"  ;
    if (arc_index == 751) return "H"  ;
    if (arc_index == 770) return "H"  ;
    if (arc_index == 779) return "H"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 797) return "E"  ;
    if (arc_index == 799) return "E"  ;
    if (arc_index == 803) return "E"  ;
    if (arc_index == 808) return "E"  ;
    if (arc_index == 809) return "W"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 812) return "E"  ;
    if (arc_index == 829) return "H"  ;
    if (arc_index == 865) return "H"  ;
    if (arc_index == 900) return "H"  ;
    if (arc_index == 902) return "H"  ;
    if (arc_index == 912) return "W"  ;
    if (arc_index == 915) return "W"  ;
    if (arc_index == 918) return "H"  ;
    if (arc_index == 924) return "W"  ;
    if (arc_index == 931) return "W"  ;
    if (arc_index == 932) return "H"  ;
    if (arc_index == 935) return "H"  ;
    if (arc_index == 938) return "W"  ;
    if (arc_index == 942) return "W"  ;
    if (arc_index == 946) return "E"  ;
    if (arc_index == 957) return "E"  ;
    if (arc_index == 978) return "W"  ;
    if (arc_index == 1010) return "W"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1029) return "E"  ;
    if (arc_index == 1032) return "E"  ;
    if (arc_index == 1063) return "H"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1179) return "W"  ;
    if (arc_index == 1190) return "W"  ;
    if (arc_index == 1191) return "W"  ;
    if (arc_index == 1192) return "W"  ;
    if (arc_index == 1193) return "W"  ;
    if (arc_index == 1197) return "W"  ;
    if (arc_index == 1202) return "W"  ;
    if (arc_index == 1205) return "W"  ;
    if (arc_index == 1208) return "W"  ;
    if (arc_index == 1209) return "W"  ;
    if (arc_index == 1216) return "H"  ;
    if (arc_index == 1220) return "H"  ;
    if (arc_index == 1231) return "H"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1292) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1437) return "W"  ;
    if (arc_index == 1465) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1499) return "W"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1533) return "W"  ;
    if (arc_index == 1538) return "E"  ;
    if (arc_index == 1539) return "E"  ;
    if (arc_index == 1563) return "E"  ;
    if (arc_index == 1637) return "E"  ;
    if (arc_index == 1642) return "E"  ;
    if (arc_index == 1644) return "E"  ;
    if (arc_index == 1659) return "W"  ;
    if (arc_index == 1719) return "E"  ;
    if (arc_index == 1723) return "E"  ;
    if (arc_index == 1726) return "E"  ;
    if (arc_index == 1735) return "E"  ;
    if (arc_index == 1740) return "E"  ;
    if (arc_index == 1743) return "E"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1789) return "E"  ;
    if (arc_index == 1790) return "E"  ;
    if (arc_index == 1795) return "E"  ;
    if (arc_index == 1835) return "E"  ;
    if (arc_index == 1865) return "H"  ;
    if (arc_index == 1921) return "H"  ;
    if (arc_index == 1929) return "E"  ;
    if (arc_index == 1935) return "E"  ;
    if (arc_index == 1937) return "E"  ;
    if (arc_index == 1972) return "E"  ;
    if (arc_index == 2002) return "E"  ;
    if (arc_index == 2007) return "E"  ;
    if (arc_index == 2013) return "E"  ;
    if (arc_index == 2014) return "W"  ;
    if (arc_index == 2015) return "W"  ;
    if (arc_index == 2020) return "H"  ;
    if (arc_index == 2021) return "W"  ;
    if (arc_index == 2035) return "W"  ;
    if (arc_index == 2040) return "W"  ;
    if (arc_index == 2054) return "W"  ;
    if (arc_index == 2153) return "H"  ;
    if (arc_index == 2161) return "H"  ;
    if (arc_index == 2162) return "H"  ;
    if (arc_index == 2165) return "W"  ;
    if (arc_index == 2173) return "W"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2226) return "E"  ;
    if (arc_index == 2234) return "E"  ;
    if (arc_index == 2248) return "H"  ;
    if (arc_index == 2275) return "H"  ;
    if (arc_index == 2283) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2374) return "H"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2423) return "W"  ;
    if (arc_index == 2438) return "W"  ;
    if (arc_index == 2452) return "W"  ;
    if (arc_index == 2469) return "W"  ;
    if (arc_index == 2485) return "H"  ;
    if (arc_index == 2526) return "H"  ;
    if (arc_index == 2527) return "W"  ;
    if (arc_index == 2535) return "W"  ;
    if (arc_index == 2555) return "H"  ;
    if (arc_index == 2580) return "E"  ;
    if (arc_index == 2589) return "E"  ;
    if (arc_index == 2590) return "E"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2672) return "E"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2730) return "H"  ;
    if (arc_index == 2733) return "H"  ;
    if (arc_index == 2746) return "H"  ;
    if (arc_index == 2765) return "H"  ;
    if (arc_index == 2793) return "H"  ;
    if (arc_index == 2812) return "E"  ;
    if (arc_index == 2868) return "E"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 7)) begin 
    if (arc_index == 23) return "H"  ;
    if (arc_index == 66) return "H"  ;
    if (arc_index == 88) return "W"  ;
    if (arc_index == 89) return "E"  ;
    if (arc_index == 90) return "E"  ;
    if (arc_index == 91) return "E"  ;
    if (arc_index == 92) return "E"  ;
    if (arc_index == 93) return "W"  ;
    if (arc_index == 94) return "E"  ;
    if (arc_index == 95) return "E"  ;
    if (arc_index == 96) return "W"  ;
    if (arc_index == 97) return "W"  ;
    if (arc_index == 98) return "W"  ;
    if (arc_index == 99) return "W"  ;
    if (arc_index == 100) return "W"  ;
    if (arc_index == 101) return "W"  ;
    if (arc_index == 102) return "W"  ;
    if (arc_index == 103) return "W"  ;
    if (arc_index == 104) return "E"  ;
    if (arc_index == 105) return "E"  ;
    if (arc_index == 106) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 108) return "W"  ;
    if (arc_index == 109) return "W"  ;
    if (arc_index == 111) return "E"  ;
    if (arc_index == 121) return "H"  ;
    if (arc_index == 126) return "H"  ;
    if (arc_index == 127) return "E"  ;
    if (arc_index == 147) return "E"  ;
    if (arc_index == 156) return "E"  ;
    if (arc_index == 166) return "H"  ;
    if (arc_index == 237) return "H"  ;
    if (arc_index == 287) return "H"  ;
    if (arc_index == 354) return "H"  ;
    if (arc_index == 365) return "H"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 393) return "E"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 401) return "E"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 415) return "E"  ;
    if (arc_index == 420) return "E"  ;
    if (arc_index == 422) return "E"  ;
    if (arc_index == 426) return "W"  ;
    if (arc_index == 428) return "W"  ;
    if (arc_index == 431) return "W"  ;
    if (arc_index == 433) return "W"  ;
    if (arc_index == 436) return "W"  ;
    if (arc_index == 437) return "W"  ;
    if (arc_index == 438) return "W"  ;
    if (arc_index == 451) return "W"  ;
    if (arc_index == 459) return "W"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 533) return "E"  ;
    if (arc_index == 542) return "H"  ;
    if (arc_index == 596) return "W"  ;
    if (arc_index == 616) return "W"  ;
    if (arc_index == 626) return "H"  ;
    if (arc_index == 643) return "H"  ;
    if (arc_index == 646) return "H"  ;
    if (arc_index == 652) return "H"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 695) return "E"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 726) return "W"  ;
    if (arc_index == 729) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 735) return "H"  ;
    if (arc_index == 742) return "H"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 759) return "E"  ;
    if (arc_index == 795) return "E"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 851) return "H"  ;
    if (arc_index == 857) return "H"  ;
    if (arc_index == 933) return "H"  ;
    if (arc_index == 940) return "H"  ;
    if (arc_index == 941) return "E"  ;
    if (arc_index == 954) return "H"  ;
    if (arc_index == 956) return "H"  ;
    if (arc_index == 970) return "E"  ;
    if (arc_index == 992) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1044) return "E"  ;
    if (arc_index == 1046) return "E"  ;
    if (arc_index == 1047) return "E"  ;
    if (arc_index == 1065) return "E"  ;
    if (arc_index == 1085) return "H"  ;
    if (arc_index == 1102) return "H"  ;
    if (arc_index == 1139) return "H"  ;
    if (arc_index == 1159) return "H"  ;
    if (arc_index == 1163) return "H"  ;
    if (arc_index == 1189) return "E"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1234) return "E"  ;
    if (arc_index == 1238) return "H"  ;
    if (arc_index == 1240) return "W"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1245) return "W"  ;
    if (arc_index == 1246) return "W"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1258) return "W"  ;
    if (arc_index == 1260) return "W"  ;
    if (arc_index == 1262) return "W"  ;
    if (arc_index == 1267) return "W"  ;
    if (arc_index == 1272) return "W"  ;
    if (arc_index == 1282) return "W"  ;
    if (arc_index == 1284) return "W"  ;
    if (arc_index == 1285) return "W"  ;
    if (arc_index == 1287) return "E"  ;
    if (arc_index == 1301) return "E"  ;
    if (arc_index == 1303) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1309) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1367) return "W"  ;
    if (arc_index == 1370) return "W"  ;
    if (arc_index == 1374) return "W"  ;
    if (arc_index == 1375) return "W"  ;
    if (arc_index == 1377) return "W"  ;
    if (arc_index == 1379) return "W"  ;
    if (arc_index == 1380) return "W"  ;
    if (arc_index == 1382) return "E"  ;
    if (arc_index == 1385) return "E"  ;
    if (arc_index == 1397) return "E"  ;
    if (arc_index == 1415) return "E"  ;
    if (arc_index == 1442) return "E"  ;
    if (arc_index == 1509) return "E"  ;
    if (arc_index == 1510) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1641) return "E"  ;
    if (arc_index == 1677) return "W"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1810) return "W"  ;
    if (arc_index == 1818) return "W"  ;
    if (arc_index == 1887) return "H"  ;
    if (arc_index == 1890) return "W"  ;
    if (arc_index == 1902) return "W"  ;
    if (arc_index == 1945) return "W"  ;
    if (arc_index == 1988) return "W"  ;
    if (arc_index == 2010) return "W"  ;
    if (arc_index == 2019) return "W"  ;
    if (arc_index == 2031) return "W"  ;
    if (arc_index == 2042) return "H"  ;
    if (arc_index == 2061) return "H"  ;
    if (arc_index == 2069) return "W"  ;
    if (arc_index == 2071) return "W"  ;
    if (arc_index == 2074) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2120) return "E"  ;
    if (arc_index == 2127) return "E"  ;
    if (arc_index == 2136) return "E"  ;
    if (arc_index == 2142) return "E"  ;
    if (arc_index == 2146) return "E"  ;
    if (arc_index == 2147) return "E"  ;
    if (arc_index == 2175) return "H"  ;
    if (arc_index == 2183) return "H"  ;
    if (arc_index == 2195) return "H"  ;
    if (arc_index == 2197) return "W"  ;
    if (arc_index == 2201) return "W"  ;
    if (arc_index == 2202) return "W"  ;
    if (arc_index == 2205) return "W"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2251) return "E"  ;
    if (arc_index == 2270) return "H"  ;
    if (arc_index == 2348) return "H"  ;
    if (arc_index == 2372) return "H"  ;
    if (arc_index == 2396) return "H"  ;
    if (arc_index == 2411) return "W"  ;
    if (arc_index == 2418) return "W"  ;
    if (arc_index == 2428) return "E"  ;
    if (arc_index == 2444) return "E"  ;
    if (arc_index == 2446) return "E"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2505) return "E"  ;
    if (arc_index == 2507) return "H"  ;
    if (arc_index == 2517) return "H"  ;
    if (arc_index == 2522) return "E"  ;
    if (arc_index == 2525) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2577) return "H"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2600) return "E"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2719) return "W"  ;
    if (arc_index == 2725) return "W"  ;
    if (arc_index == 2752) return "H"  ;
    if (arc_index == 2837) return "H"  ;
    if (arc_index == 2907) return "H"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 5)) begin 
    if (arc_index == 23) return "E"  ;
    if (arc_index == 37) return "E"  ;
    if (arc_index == 45) return "H"  ;
    if (arc_index == 66) return "E"  ;
    if (arc_index == 88) return "H"  ;
    if (arc_index == 93) return "W"  ;
    if (arc_index == 96) return "W"  ;
    if (arc_index == 99) return "W"  ;
    if (arc_index == 102) return "W"  ;
    if (arc_index == 110) return "W"  ;
    if (arc_index == 111) return "E"  ;
    if (arc_index == 112) return "W"  ;
    if (arc_index == 113) return "W"  ;
    if (arc_index == 114) return "W"  ;
    if (arc_index == 115) return "W"  ;
    if (arc_index == 116) return "W"  ;
    if (arc_index == 117) return "W"  ;
    if (arc_index == 118) return "W"  ;
    if (arc_index == 119) return "W"  ;
    if (arc_index == 120) return "W"  ;
    if (arc_index == 121) return "E"  ;
    if (arc_index == 122) return "E"  ;
    if (arc_index == 123) return "E"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 125) return "E"  ;
    if (arc_index == 126) return "E"  ;
    if (arc_index == 127) return "E"  ;
    if (arc_index == 128) return "E"  ;
    if (arc_index == 129) return "E"  ;
    if (arc_index == 130) return "E"  ;
    if (arc_index == 131) return "E"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 137) return "E"  ;
    if (arc_index == 143) return "H"  ;
    if (arc_index == 149) return "H"  ;
    if (arc_index == 163) return "W"  ;
    if (arc_index == 165) return "W"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 188) return "H"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 331) return "W"  ;
    if (arc_index == 345) return "W"  ;
    if (arc_index == 358) return "W"  ;
    if (arc_index == 371) return "W"  ;
    if (arc_index == 374) return "W"  ;
    if (arc_index == 376) return "E"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 385) return "E"  ;
    if (arc_index == 387) return "H"  ;
    if (arc_index == 393) return "E"  ;
    if (arc_index == 397) return "W"  ;
    if (arc_index == 399) return "W"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 401) return "E"  ;
    if (arc_index == 402) return "E"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 404) return "E"  ;
    if (arc_index == 405) return "W"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 408) return "E"  ;
    if (arc_index == 410) return "W"  ;
    if (arc_index == 412) return "W"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 414) return "E"  ;
    if (arc_index == 415) return "E"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 451) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 474) return "E"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 564) return "H"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 640) return "E"  ;
    if (arc_index == 641) return "W"  ;
    if (arc_index == 644) return "W"  ;
    if (arc_index == 645) return "W"  ;
    if (arc_index == 648) return "H"  ;
    if (arc_index == 650) return "H"  ;
    if (arc_index == 651) return "W"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 677) return "E"  ;
    if (arc_index == 752) return "E"  ;
    if (arc_index == 757) return "H"  ;
    if (arc_index == 795) return "E"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 850) return "W"  ;
    if (arc_index == 862) return "W"  ;
    if (arc_index == 873) return "H"  ;
    if (arc_index == 874) return "H"  ;
    if (arc_index == 879) return "H"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 915) return "E"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 940) return "E"  ;
    if (arc_index == 941) return "E"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 962) return "H"  ;
    if (arc_index == 968) return "H"  ;
    if (arc_index == 970) return "E"  ;
    if (arc_index == 976) return "H"  ;
    if (arc_index == 984) return "H"  ;
    if (arc_index == 989) return "H"  ;
    if (arc_index == 991) return "H"  ;
    if (arc_index == 1001) return "H"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1041) return "W"  ;
    if (arc_index == 1059) return "W"  ;
    if (arc_index == 1107) return "H"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1240) return "W"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1245) return "W"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1260) return "H"  ;
    if (arc_index == 1262) return "H"  ;
    if (arc_index == 1267) return "W"  ;
    if (arc_index == 1282) return "W"  ;
    if (arc_index == 1289) return "W"  ;
    if (arc_index == 1295) return "W"  ;
    if (arc_index == 1303) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1393) return "W"  ;
    if (arc_index == 1431) return "W"  ;
    if (arc_index == 1447) return "W"  ;
    if (arc_index == 1474) return "W"  ;
    if (arc_index == 1498) return "W"  ;
    if (arc_index == 1499) return "W"  ;
    if (arc_index == 1500) return "W"  ;
    if (arc_index == 1504) return "E"  ;
    if (arc_index == 1506) return "E"  ;
    if (arc_index == 1507) return "E"  ;
    if (arc_index == 1508) return "E"  ;
    if (arc_index == 1509) return "E"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1514) return "W"  ;
    if (arc_index == 1515) return "W"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1529) return "W"  ;
    if (arc_index == 1546) return "W"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1592) return "W"  ;
    if (arc_index == 1621) return "E"  ;
    if (arc_index == 1635) return "E"  ;
    if (arc_index == 1677) return "W"  ;
    if (arc_index == 1687) return "W"  ;
    if (arc_index == 1710) return "W"  ;
    if (arc_index == 1723) return "W"  ;
    if (arc_index == 1764) return "W"  ;
    if (arc_index == 1773) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1855) return "W"  ;
    if (arc_index == 1872) return "W"  ;
    if (arc_index == 1878) return "W"  ;
    if (arc_index == 1890) return "W"  ;
    if (arc_index == 1902) return "E"  ;
    if (arc_index == 1909) return "H"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2061) return "E"  ;
    if (arc_index == 2064) return "H"  ;
    if (arc_index == 2069) return "W"  ;
    if (arc_index == 2071) return "W"  ;
    if (arc_index == 2074) return "W"  ;
    if (arc_index == 2112) return "W"  ;
    if (arc_index == 2119) return "W"  ;
    if (arc_index == 2135) return "E"  ;
    if (arc_index == 2136) return "E"  ;
    if (arc_index == 2142) return "E"  ;
    if (arc_index == 2143) return "E"  ;
    if (arc_index == 2146) return "E"  ;
    if (arc_index == 2147) return "E"  ;
    if (arc_index == 2175) return "E"  ;
    if (arc_index == 2197) return "H"  ;
    if (arc_index == 2202) return "H"  ;
    if (arc_index == 2204) return "H"  ;
    if (arc_index == 2205) return "H"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2212) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2246) return "W"  ;
    if (arc_index == 2259) return "W"  ;
    if (arc_index == 2292) return "H"  ;
    if (arc_index == 2350) return "H"  ;
    if (arc_index == 2362) return "H"  ;
    if (arc_index == 2411) return "W"  ;
    if (arc_index == 2418) return "H"  ;
    if (arc_index == 2437) return "E"  ;
    if (arc_index == 2446) return "E"  ;
    if (arc_index == 2449) return "E"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2483) return "E"  ;
    if (arc_index == 2491) return "E"  ;
    if (arc_index == 2493) return "E"  ;
    if (arc_index == 2512) return "E"  ;
    if (arc_index == 2517) return "E"  ;
    if (arc_index == 2522) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2525) return "E"  ;
    if (arc_index == 2528) return "E"  ;
    if (arc_index == 2529) return "H"  ;
    if (arc_index == 2592) return "E"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2599) return "H"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2704) return "E"  ;
    if (arc_index == 2719) return "W"  ;
    if (arc_index == 2733) return "E"  ;
    if (arc_index == 2774) return "H"  ;
    if (arc_index == 2815) return "H"  ;
    if (arc_index == 2885) return "H"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 4)) begin 
    if (arc_index == 40) return "W"  ;
    if (arc_index == 67) return "H"  ;
    if (arc_index == 110) return "H"  ;
    if (arc_index == 132) return "H"  ;
    if (arc_index == 133) return "H"  ;
    if (arc_index == 134) return "E"  ;
    if (arc_index == 135) return "E"  ;
    if (arc_index == 136) return "E"  ;
    if (arc_index == 137) return "E"  ;
    if (arc_index == 138) return "E"  ;
    if (arc_index == 139) return "E"  ;
    if (arc_index == 140) return "E"  ;
    if (arc_index == 141) return "W"  ;
    if (arc_index == 142) return "W"  ;
    if (arc_index == 143) return "E"  ;
    if (arc_index == 144) return "W"  ;
    if (arc_index == 145) return "W"  ;
    if (arc_index == 146) return "E"  ;
    if (arc_index == 147) return "E"  ;
    if (arc_index == 148) return "E"  ;
    if (arc_index == 149) return "E"  ;
    if (arc_index == 150) return "E"  ;
    if (arc_index == 151) return "W"  ;
    if (arc_index == 152) return "W"  ;
    if (arc_index == 153) return "W"  ;
    if (arc_index == 165) return "H"  ;
    if (arc_index == 210) return "H"  ;
    if (arc_index == 223) return "W"  ;
    if (arc_index == 398) return "W"  ;
    if (arc_index == 407) return "W"  ;
    if (arc_index == 409) return "H"  ;
    if (arc_index == 411) return "W"  ;
    if (arc_index == 417) return "W"  ;
    if (arc_index == 586) return "H"  ;
    if (arc_index == 595) return "W"  ;
    if (arc_index == 660) return "E"  ;
    if (arc_index == 661) return "E"  ;
    if (arc_index == 665) return "E"  ;
    if (arc_index == 669) return "E"  ;
    if (arc_index == 670) return "H"  ;
    if (arc_index == 671) return "E"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 673) return "E"  ;
    if (arc_index == 677) return "E"  ;
    if (arc_index == 680) return "E"  ;
    if (arc_index == 727) return "E"  ;
    if (arc_index == 732) return "E"  ;
    if (arc_index == 738) return "W"  ;
    if (arc_index == 779) return "H"  ;
    if (arc_index == 804) return "E"  ;
    if (arc_index == 858) return "E"  ;
    if (arc_index == 859) return "W"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 870) return "W"  ;
    if (arc_index == 875) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 895) return "H"  ;
    if (arc_index == 934) return "E"  ;
    if (arc_index == 936) return "E"  ;
    if (arc_index == 984) return "H"  ;
    if (arc_index == 998) return "H"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1114) return "W"  ;
    if (arc_index == 1129) return "H"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1171) return "W"  ;
    if (arc_index == 1258) return "W"  ;
    if (arc_index == 1282) return "H"  ;
    if (arc_index == 1307) return "W"  ;
    if (arc_index == 1378) return "W"  ;
    if (arc_index == 1384) return "W"  ;
    if (arc_index == 1512) return "W"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1565) return "W"  ;
    if (arc_index == 1724) return "E"  ;
    if (arc_index == 1810) return "W"  ;
    if (arc_index == 1931) return "H"  ;
    if (arc_index == 1980) return "W"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2005) return "E"  ;
    if (arc_index == 2008) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2011) return "E"  ;
    if (arc_index == 2016) return "E"  ;
    if (arc_index == 2018) return "E"  ;
    if (arc_index == 2019) return "E"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2086) return "H"  ;
    if (arc_index == 2219) return "H"  ;
    if (arc_index == 2227) return "H"  ;
    if (arc_index == 2230) return "E"  ;
    if (arc_index == 2279) return "W"  ;
    if (arc_index == 2314) return "H"  ;
    if (arc_index == 2440) return "H"  ;
    if (arc_index == 2459) return "W"  ;
    if (arc_index == 2514) return "E"  ;
    if (arc_index == 2551) return "H"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2621) return "H"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2796) return "H"  ;
    if (arc_index == 2812) return "E"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 8)) begin 
    if (arc_index == 11) return "E"  ;
    if (arc_index == 17) return "E"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 89) return "H"  ;
    if (arc_index == 109) return "E"  ;
    if (arc_index == 132) return "H"  ;
    if (arc_index == 154) return "H"  ;
    if (arc_index == 155) return "H"  ;
    if (arc_index == 156) return "H"  ;
    if (arc_index == 157) return "H"  ;
    if (arc_index == 158) return "W"  ;
    if (arc_index == 159) return "W"  ;
    if (arc_index == 160) return "W"  ;
    if (arc_index == 161) return "W"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 163) return "W"  ;
    if (arc_index == 164) return "W"  ;
    if (arc_index == 165) return "W"  ;
    if (arc_index == 166) return "W"  ;
    if (arc_index == 167) return "W"  ;
    if (arc_index == 168) return "E"  ;
    if (arc_index == 169) return "E"  ;
    if (arc_index == 170) return "E"  ;
    if (arc_index == 171) return "E"  ;
    if (arc_index == 172) return "E"  ;
    if (arc_index == 173) return "E"  ;
    if (arc_index == 174) return "E"  ;
    if (arc_index == 175) return "E"  ;
    if (arc_index == 177) return "E"  ;
    if (arc_index == 187) return "H"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 199) return "W"  ;
    if (arc_index == 213) return "E"  ;
    if (arc_index == 220) return "E"  ;
    if (arc_index == 228) return "E"  ;
    if (arc_index == 231) return "E"  ;
    if (arc_index == 232) return "H"  ;
    if (arc_index == 242) return "H"  ;
    if (arc_index == 249) return "H"  ;
    if (arc_index == 250) return "H"  ;
    if (arc_index == 252) return "H"  ;
    if (arc_index == 253) return "H"  ;
    if (arc_index == 260) return "H"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 275) return "W"  ;
    if (arc_index == 276) return "W"  ;
    if (arc_index == 278) return "W"  ;
    if (arc_index == 281) return "W"  ;
    if (arc_index == 288) return "W"  ;
    if (arc_index == 308) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 327) return "W"  ;
    if (arc_index == 347) return "W"  ;
    if (arc_index == 354) return "W"  ;
    if (arc_index == 377) return "W"  ;
    if (arc_index == 386) return "W"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 420) return "E"  ;
    if (arc_index == 431) return "H"  ;
    if (arc_index == 502) return "H"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 528) return "E"  ;
    if (arc_index == 547) return "E"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 608) return "H"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 613) return "W"  ;
    if (arc_index == 619) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 643) return "W"  ;
    if (arc_index == 660) return "W"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 689) return "E"  ;
    if (arc_index == 692) return "H"  ;
    if (arc_index == 695) return "H"  ;
    if (arc_index == 700) return "H"  ;
    if (arc_index == 702) return "H"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 718) return "W"  ;
    if (arc_index == 721) return "W"  ;
    if (arc_index == 730) return "W"  ;
    if (arc_index == 758) return "W"  ;
    if (arc_index == 801) return "H"  ;
    if (arc_index == 833) return "H"  ;
    if (arc_index == 841) return "H"  ;
    if (arc_index == 882) return "E"  ;
    if (arc_index == 883) return "E"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 917) return "H"  ;
    if (arc_index == 929) return "H"  ;
    if (arc_index == 1006) return "H"  ;
    if (arc_index == 1020) return "H"  ;
    if (arc_index == 1040) return "H"  ;
    if (arc_index == 1050) return "W"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1103) return "E"  ;
    if (arc_index == 1118) return "E"  ;
    if (arc_index == 1136) return "E"  ;
    if (arc_index == 1144) return "E"  ;
    if (arc_index == 1145) return "E"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1148) return "W"  ;
    if (arc_index == 1149) return "W"  ;
    if (arc_index == 1150) return "W"  ;
    if (arc_index == 1151) return "H"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1161) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1164) return "W"  ;
    if (arc_index == 1165) return "W"  ;
    if (arc_index == 1177) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1236) return "E"  ;
    if (arc_index == 1239) return "E"  ;
    if (arc_index == 1251) return "E"  ;
    if (arc_index == 1257) return "W"  ;
    if (arc_index == 1259) return "W"  ;
    if (arc_index == 1263) return "W"  ;
    if (arc_index == 1304) return "H"  ;
    if (arc_index == 1329) return "H"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1341) return "W"  ;
    if (arc_index == 1344) return "W"  ;
    if (arc_index == 1394) return "E"  ;
    if (arc_index == 1398) return "E"  ;
    if (arc_index == 1399) return "E"  ;
    if (arc_index == 1410) return "E"  ;
    if (arc_index == 1414) return "E"  ;
    if (arc_index == 1426) return "E"  ;
    if (arc_index == 1445) return "E"  ;
    if (arc_index == 1460) return "E"  ;
    if (arc_index == 1474) return "E"  ;
    if (arc_index == 1475) return "E"  ;
    if (arc_index == 1479) return "E"  ;
    if (arc_index == 1480) return "E"  ;
    if (arc_index == 1487) return "E"  ;
    if (arc_index == 1488) return "E"  ;
    if (arc_index == 1489) return "E"  ;
    if (arc_index == 1490) return "E"  ;
    if (arc_index == 1501) return "E"  ;
    if (arc_index == 1507) return "E"  ;
    if (arc_index == 1515) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1544) return "E"  ;
    if (arc_index == 1554) return "W"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1610) return "E"  ;
    if (arc_index == 1613) return "E"  ;
    if (arc_index == 1619) return "E"  ;
    if (arc_index == 1654) return "E"  ;
    if (arc_index == 1679) return "E"  ;
    if (arc_index == 1680) return "E"  ;
    if (arc_index == 1685) return "E"  ;
    if (arc_index == 1688) return "E"  ;
    if (arc_index == 1705) return "E"  ;
    if (arc_index == 1708) return "E"  ;
    if (arc_index == 1736) return "E"  ;
    if (arc_index == 1763) return "E"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1787) return "E"  ;
    if (arc_index == 1791) return "E"  ;
    if (arc_index == 1792) return "E"  ;
    if (arc_index == 1797) return "E"  ;
    if (arc_index == 1805) return "E"  ;
    if (arc_index == 1806) return "E"  ;
    if (arc_index == 1809) return "E"  ;
    if (arc_index == 1817) return "E"  ;
    if (arc_index == 1825) return "E"  ;
    if (arc_index == 1847) return "E"  ;
    if (arc_index == 1858) return "E"  ;
    if (arc_index == 1867) return "E"  ;
    if (arc_index == 1869) return "E"  ;
    if (arc_index == 1882) return "W"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1917) return "E"  ;
    if (arc_index == 1953) return "H"  ;
    if (arc_index == 1964) return "H"  ;
    if (arc_index == 1995) return "H"  ;
    if (arc_index == 2012) return "H"  ;
    if (arc_index == 2072) return "H"  ;
    if (arc_index == 2081) return "W"  ;
    if (arc_index == 2098) return "W"  ;
    if (arc_index == 2106) return "W"  ;
    if (arc_index == 2108) return "H"  ;
    if (arc_index == 2121) return "H"  ;
    if (arc_index == 2160) return "H"  ;
    if (arc_index == 2214) return "H"  ;
    if (arc_index == 2237) return "H"  ;
    if (arc_index == 2241) return "H"  ;
    if (arc_index == 2249) return "H"  ;
    if (arc_index == 2294) return "E"  ;
    if (arc_index == 2303) return "E"  ;
    if (arc_index == 2307) return "E"  ;
    if (arc_index == 2313) return "W"  ;
    if (arc_index == 2329) return "W"  ;
    if (arc_index == 2336) return "H"  ;
    if (arc_index == 2338) return "H"  ;
    if (arc_index == 2344) return "H"  ;
    if (arc_index == 2352) return "H"  ;
    if (arc_index == 2355) return "H"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2359) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2363) return "W"  ;
    if (arc_index == 2364) return "W"  ;
    if (arc_index == 2366) return "W"  ;
    if (arc_index == 2367) return "W"  ;
    if (arc_index == 2368) return "W"  ;
    if (arc_index == 2369) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2372) return "W"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2375) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2432) return "E"  ;
    if (arc_index == 2462) return "H"  ;
    if (arc_index == 2468) return "H"  ;
    if (arc_index == 2470) return "H"  ;
    if (arc_index == 2476) return "H"  ;
    if (arc_index == 2482) return "H"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2573) return "H"  ;
    if (arc_index == 2600) return "H"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2620) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2627) return "W"  ;
    if (arc_index == 2643) return "H"  ;
    if (arc_index == 2645) return "H"  ;
    if (arc_index == 2661) return "H"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2753) return "W"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2818) return "H"  ;
    if (arc_index == 2822) return "H"  ;
    if (arc_index == 2831) return "H"  ;
    if (arc_index == 2848) return "H"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2892) return "E"  ;
    if (arc_index == 2912) return "W"  ;
    if (arc_index == 2915) return "W"  ;
    if (arc_index == 2919) return "W"  ;
    if (arc_index == 2922) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 10)) begin 
    if (arc_index == 62) return "E"  ;
    if (arc_index == 104) return "E"  ;
    if (arc_index == 111) return "H"  ;
    if (arc_index == 146) return "E"  ;
    if (arc_index == 154) return "H"  ;
    if (arc_index == 176) return "W"  ;
    if (arc_index == 177) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 179) return "W"  ;
    if (arc_index == 180) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 182) return "W"  ;
    if (arc_index == 183) return "W"  ;
    if (arc_index == 184) return "W"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 187) return "W"  ;
    if (arc_index == 188) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 191) return "W"  ;
    if (arc_index == 192) return "W"  ;
    if (arc_index == 193) return "W"  ;
    if (arc_index == 194) return "W"  ;
    if (arc_index == 195) return "E"  ;
    if (arc_index == 196) return "E"  ;
    if (arc_index == 197) return "E"  ;
    if (arc_index == 203) return "E"  ;
    if (arc_index == 209) return "H"  ;
    if (arc_index == 254) return "H"  ;
    if (arc_index == 283) return "H"  ;
    if (arc_index == 289) return "H"  ;
    if (arc_index == 290) return "E"  ;
    if (arc_index == 291) return "E"  ;
    if (arc_index == 292) return "E"  ;
    if (arc_index == 304) return "W"  ;
    if (arc_index == 370) return "W"  ;
    if (arc_index == 453) return "H"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 614) return "E"  ;
    if (arc_index == 615) return "E"  ;
    if (arc_index == 630) return "H"  ;
    if (arc_index == 646) return "H"  ;
    if (arc_index == 672) return "H"  ;
    if (arc_index == 685) return "H"  ;
    if (arc_index == 714) return "H"  ;
    if (arc_index == 723) return "H"  ;
    if (arc_index == 740) return "H"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 818) return "E"  ;
    if (arc_index == 823) return "H"  ;
    if (arc_index == 939) return "H"  ;
    if (arc_index == 969) return "E"  ;
    if (arc_index == 1028) return "H"  ;
    if (arc_index == 1037) return "H"  ;
    if (arc_index == 1042) return "H"  ;
    if (arc_index == 1053) return "H"  ;
    if (arc_index == 1057) return "H"  ;
    if (arc_index == 1067) return "E"  ;
    if (arc_index == 1100) return "E"  ;
    if (arc_index == 1112) return "E"  ;
    if (arc_index == 1122) return "E"  ;
    if (arc_index == 1124) return "W"  ;
    if (arc_index == 1127) return "W"  ;
    if (arc_index == 1128) return "W"  ;
    if (arc_index == 1130) return "W"  ;
    if (arc_index == 1132) return "W"  ;
    if (arc_index == 1133) return "W"  ;
    if (arc_index == 1134) return "W"  ;
    if (arc_index == 1136) return "W"  ;
    if (arc_index == 1138) return "W"  ;
    if (arc_index == 1140) return "W"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1142) return "W"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1155) return "W"  ;
    if (arc_index == 1173) return "H"  ;
    if (arc_index == 1241) return "H"  ;
    if (arc_index == 1249) return "H"  ;
    if (arc_index == 1324) return "H"  ;
    if (arc_index == 1326) return "H"  ;
    if (arc_index == 1399) return "H"  ;
    if (arc_index == 1450) return "H"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1561) return "W"  ;
    if (arc_index == 1567) return "W"  ;
    if (arc_index == 1570) return "W"  ;
    if (arc_index == 1577) return "W"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1583) return "W"  ;
    if (arc_index == 1595) return "W"  ;
    if (arc_index == 1660) return "W"  ;
    if (arc_index == 1769) return "W"  ;
    if (arc_index == 1797) return "E"  ;
    if (arc_index == 1806) return "E"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1886) return "E"  ;
    if (arc_index == 1975) return "H"  ;
    if (arc_index == 2068) return "H"  ;
    if (arc_index == 2070) return "H"  ;
    if (arc_index == 2072) return "W"  ;
    if (arc_index == 2073) return "W"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2077) return "W"  ;
    if (arc_index == 2078) return "W"  ;
    if (arc_index == 2079) return "W"  ;
    if (arc_index == 2081) return "W"  ;
    if (arc_index == 2083) return "W"  ;
    if (arc_index == 2085) return "W"  ;
    if (arc_index == 2087) return "W"  ;
    if (arc_index == 2088) return "W"  ;
    if (arc_index == 2089) return "W"  ;
    if (arc_index == 2100) return "W"  ;
    if (arc_index == 2101) return "W"  ;
    if (arc_index == 2130) return "H"  ;
    if (arc_index == 2133) return "E"  ;
    if (arc_index == 2178) return "E"  ;
    if (arc_index == 2180) return "W"  ;
    if (arc_index == 2184) return "W"  ;
    if (arc_index == 2195) return "W"  ;
    if (arc_index == 2197) return "W"  ;
    if (arc_index == 2208) return "W"  ;
    if (arc_index == 2211) return "W"  ;
    if (arc_index == 2263) return "H"  ;
    if (arc_index == 2271) return "H"  ;
    if (arc_index == 2311) return "H"  ;
    if (arc_index == 2345) return "H"  ;
    if (arc_index == 2358) return "H"  ;
    if (arc_index == 2382) return "H"  ;
    if (arc_index == 2388) return "W"  ;
    if (arc_index == 2414) return "W"  ;
    if (arc_index == 2444) return "W"  ;
    if (arc_index == 2455) return "W"  ;
    if (arc_index == 2484) return "H"  ;
    if (arc_index == 2595) return "H"  ;
    if (arc_index == 2606) return "H"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2665) return "H"  ;
    if (arc_index == 2712) return "H"  ;
    if (arc_index == 2715) return "H"  ;
    if (arc_index == 2719) return "W"  ;
    if (arc_index == 2725) return "W"  ;
    if (arc_index == 2831) return "W"  ;
    if (arc_index == 2840) return "H"  ;
    if (arc_index == 2920) return "H"  ;
    if (arc_index == 2921) return "H"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 7)) begin 
    if (arc_index == 9) return "H"  ;
    if (arc_index == 16) return "H"  ;
    if (arc_index == 43) return "H"  ;
    if (arc_index == 92) return "W"  ;
    if (arc_index == 95) return "W"  ;
    if (arc_index == 125) return "W"  ;
    if (arc_index == 133) return "H"  ;
    if (arc_index == 176) return "H"  ;
    if (arc_index == 189) return "H"  ;
    if (arc_index == 198) return "H"  ;
    if (arc_index == 199) return "E"  ;
    if (arc_index == 200) return "W"  ;
    if (arc_index == 201) return "W"  ;
    if (arc_index == 202) return "W"  ;
    if (arc_index == 203) return "E"  ;
    if (arc_index == 204) return "W"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 206) return "W"  ;
    if (arc_index == 207) return "W"  ;
    if (arc_index == 208) return "E"  ;
    if (arc_index == 209) return "E"  ;
    if (arc_index == 210) return "E"  ;
    if (arc_index == 211) return "W"  ;
    if (arc_index == 212) return "W"  ;
    if (arc_index == 213) return "E"  ;
    if (arc_index == 214) return "E"  ;
    if (arc_index == 215) return "E"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 217) return "W"  ;
    if (arc_index == 218) return "W"  ;
    if (arc_index == 219) return "W"  ;
    if (arc_index == 228) return "W"  ;
    if (arc_index == 231) return "H"  ;
    if (arc_index == 244) return "W"  ;
    if (arc_index == 261) return "W"  ;
    if (arc_index == 276) return "H"  ;
    if (arc_index == 281) return "H"  ;
    if (arc_index == 288) return "H"  ;
    if (arc_index == 300) return "H"  ;
    if (arc_index == 311) return "W"  ;
    if (arc_index == 312) return "W"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 323) return "W"  ;
    if (arc_index == 325) return "W"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 329) return "W"  ;
    if (arc_index == 359) return "W"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 475) return "H"  ;
    if (arc_index == 512) return "H"  ;
    if (arc_index == 519) return "H"  ;
    if (arc_index == 554) return "H"  ;
    if (arc_index == 557) return "H"  ;
    if (arc_index == 561) return "H"  ;
    if (arc_index == 564) return "H"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 601) return "W"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 634) return "W"  ;
    if (arc_index == 652) return "H"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 686) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 688) return "W"  ;
    if (arc_index == 690) return "W"  ;
    if (arc_index == 691) return "W"  ;
    if (arc_index == 693) return "W"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 698) return "W"  ;
    if (arc_index == 699) return "W"  ;
    if (arc_index == 710) return "W"  ;
    if (arc_index == 719) return "W"  ;
    if (arc_index == 736) return "H"  ;
    if (arc_index == 749) return "H"  ;
    if (arc_index == 758) return "H"  ;
    if (arc_index == 760) return "E"  ;
    if (arc_index == 762) return "E"  ;
    if (arc_index == 814) return "W"  ;
    if (arc_index == 827) return "W"  ;
    if (arc_index == 841) return "W"  ;
    if (arc_index == 842) return "E"  ;
    if (arc_index == 844) return "E"  ;
    if (arc_index == 845) return "H"  ;
    if (arc_index == 846) return "E"  ;
    if (arc_index == 847) return "E"  ;
    if (arc_index == 856) return "E"  ;
    if (arc_index == 892) return "E"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 961) return "H"  ;
    if (arc_index == 1004) return "H"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1050) return "H"  ;
    if (arc_index == 1064) return "H"  ;
    if (arc_index == 1088) return "H"  ;
    if (arc_index == 1108) return "H"  ;
    if (arc_index == 1161) return "H"  ;
    if (arc_index == 1174) return "E"  ;
    if (arc_index == 1195) return "H"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1313) return "E"  ;
    if (arc_index == 1316) return "E"  ;
    if (arc_index == 1321) return "W"  ;
    if (arc_index == 1348) return "H"  ;
    if (arc_index == 1374) return "W"  ;
    if (arc_index == 1379) return "E"  ;
    if (arc_index == 1399) return "E"  ;
    if (arc_index == 1404) return "E"  ;
    if (arc_index == 1409) return "E"  ;
    if (arc_index == 1414) return "E"  ;
    if (arc_index == 1427) return "E"  ;
    if (arc_index == 1449) return "E"  ;
    if (arc_index == 1460) return "E"  ;
    if (arc_index == 1476) return "W"  ;
    if (arc_index == 1486) return "W"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1544) return "E"  ;
    if (arc_index == 1558) return "W"  ;
    if (arc_index == 1624) return "W"  ;
    if (arc_index == 1670) return "W"  ;
    if (arc_index == 1688) return "W"  ;
    if (arc_index == 1714) return "E"  ;
    if (arc_index == 1739) return "E"  ;
    if (arc_index == 1764) return "E"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1793) return "E"  ;
    if (arc_index == 1816) return "W"  ;
    if (arc_index == 1828) return "W"  ;
    if (arc_index == 1832) return "E"  ;
    if (arc_index == 1851) return "E"  ;
    if (arc_index == 1895) return "E"  ;
    if (arc_index == 1997) return "H"  ;
    if (arc_index == 2093) return "W"  ;
    if (arc_index == 2095) return "W"  ;
    if (arc_index == 2097) return "W"  ;
    if (arc_index == 2103) return "W"  ;
    if (arc_index == 2104) return "W"  ;
    if (arc_index == 2123) return "E"  ;
    if (arc_index == 2152) return "H"  ;
    if (arc_index == 2168) return "H"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2215) return "W"  ;
    if (arc_index == 2262) return "E"  ;
    if (arc_index == 2266) return "E"  ;
    if (arc_index == 2285) return "H"  ;
    if (arc_index == 2288) return "H"  ;
    if (arc_index == 2292) return "H"  ;
    if (arc_index == 2293) return "H"  ;
    if (arc_index == 2294) return "H"  ;
    if (arc_index == 2295) return "E"  ;
    if (arc_index == 2296) return "E"  ;
    if (arc_index == 2299) return "E"  ;
    if (arc_index == 2302) return "W"  ;
    if (arc_index == 2303) return "W"  ;
    if (arc_index == 2306) return "W"  ;
    if (arc_index == 2307) return "W"  ;
    if (arc_index == 2308) return "W"  ;
    if (arc_index == 2309) return "W"  ;
    if (arc_index == 2321) return "W"  ;
    if (arc_index == 2335) return "W"  ;
    if (arc_index == 2346) return "W"  ;
    if (arc_index == 2366) return "W"  ;
    if (arc_index == 2380) return "H"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2467) return "E"  ;
    if (arc_index == 2471) return "E"  ;
    if (arc_index == 2476) return "E"  ;
    if (arc_index == 2481) return "E"  ;
    if (arc_index == 2482) return "E"  ;
    if (arc_index == 2503) return "E"  ;
    if (arc_index == 2504) return "E"  ;
    if (arc_index == 2506) return "H"  ;
    if (arc_index == 2538) return "H"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2603) return "W"  ;
    if (arc_index == 2605) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2608) return "W"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2617) return "H"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2635) return "W"  ;
    if (arc_index == 2637) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2687) return "H"  ;
    if (arc_index == 2757) return "E"  ;
    if (arc_index == 2769) return "E"  ;
    if (arc_index == 2776) return "E"  ;
    if (arc_index == 2777) return "E"  ;
    if (arc_index == 2786) return "E"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2816) return "E"  ;
    if (arc_index == 2826) return "E"  ;
    if (arc_index == 2829) return "E"  ;
    if (arc_index == 2832) return "W"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2862) return "H"  ;
    if (arc_index == 2864) return "E"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2923) return "W"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 8)) begin 
    if (arc_index == 21) return "E"  ;
    if (arc_index == 24) return "E"  ;
    if (arc_index == 53) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 57) return "E"  ;
    if (arc_index == 62) return "E"  ;
    if (arc_index == 89) return "E"  ;
    if (arc_index == 91) return "E"  ;
    if (arc_index == 109) return "E"  ;
    if (arc_index == 118) return "E"  ;
    if (arc_index == 119) return "E"  ;
    if (arc_index == 154) return "E"  ;
    if (arc_index == 155) return "H"  ;
    if (arc_index == 163) return "H"  ;
    if (arc_index == 166) return "H"  ;
    if (arc_index == 171) return "H"  ;
    if (arc_index == 183) return "H"  ;
    if (arc_index == 187) return "H"  ;
    if (arc_index == 192) return "W"  ;
    if (arc_index == 198) return "H"  ;
    if (arc_index == 219) return "H"  ;
    if (arc_index == 220) return "H"  ;
    if (arc_index == 221) return "E"  ;
    if (arc_index == 222) return "W"  ;
    if (arc_index == 223) return "W"  ;
    if (arc_index == 224) return "W"  ;
    if (arc_index == 225) return "W"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 227) return "W"  ;
    if (arc_index == 228) return "W"  ;
    if (arc_index == 229) return "W"  ;
    if (arc_index == 230) return "W"  ;
    if (arc_index == 231) return "W"  ;
    if (arc_index == 232) return "W"  ;
    if (arc_index == 233) return "W"  ;
    if (arc_index == 234) return "E"  ;
    if (arc_index == 235) return "E"  ;
    if (arc_index == 236) return "E"  ;
    if (arc_index == 237) return "E"  ;
    if (arc_index == 238) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 240) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 249) return "E"  ;
    if (arc_index == 252) return "E"  ;
    if (arc_index == 253) return "H"  ;
    if (arc_index == 260) return "H"  ;
    if (arc_index == 271) return "H"  ;
    if (arc_index == 279) return "H"  ;
    if (arc_index == 282) return "H"  ;
    if (arc_index == 283) return "E"  ;
    if (arc_index == 298) return "H"  ;
    if (arc_index == 299) return "W"  ;
    if (arc_index == 303) return "W"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 339) return "W"  ;
    if (arc_index == 341) return "W"  ;
    if (arc_index == 348) return "E"  ;
    if (arc_index == 364) return "E"  ;
    if (arc_index == 402) return "E"  ;
    if (arc_index == 420) return "E"  ;
    if (arc_index == 463) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 497) return "H"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 530) return "W"  ;
    if (arc_index == 531) return "W"  ;
    if (arc_index == 532) return "W"  ;
    if (arc_index == 533) return "W"  ;
    if (arc_index == 535) return "W"  ;
    if (arc_index == 537) return "W"  ;
    if (arc_index == 538) return "W"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 540) return "W"  ;
    if (arc_index == 542) return "W"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 547) return "W"  ;
    if (arc_index == 548) return "W"  ;
    if (arc_index == 554) return "W"  ;
    if (arc_index == 561) return "E"  ;
    if (arc_index == 596) return "E"  ;
    if (arc_index == 599) return "W"  ;
    if (arc_index == 616) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 636) return "W"  ;
    if (arc_index == 639) return "E"  ;
    if (arc_index == 660) return "E"  ;
    if (arc_index == 674) return "H"  ;
    if (arc_index == 704) return "H"  ;
    if (arc_index == 730) return "H"  ;
    if (arc_index == 736) return "H"  ;
    if (arc_index == 758) return "H"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 817) return "E"  ;
    if (arc_index == 867) return "H"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 982) return "E"  ;
    if (arc_index == 983) return "H"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1040) return "E"  ;
    if (arc_index == 1052) return "E"  ;
    if (arc_index == 1053) return "W"  ;
    if (arc_index == 1072) return "H"  ;
    if (arc_index == 1073) return "H"  ;
    if (arc_index == 1086) return "H"  ;
    if (arc_index == 1112) return "E"  ;
    if (arc_index == 1124) return "W"  ;
    if (arc_index == 1127) return "W"  ;
    if (arc_index == 1134) return "W"  ;
    if (arc_index == 1140) return "W"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1175) return "E"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1217) return "H"  ;
    if (arc_index == 1227) return "H"  ;
    if (arc_index == 1235) return "H"  ;
    if (arc_index == 1236) return "H"  ;
    if (arc_index == 1239) return "H"  ;
    if (arc_index == 1255) return "H"  ;
    if (arc_index == 1257) return "H"  ;
    if (arc_index == 1259) return "H"  ;
    if (arc_index == 1261) return "H"  ;
    if (arc_index == 1263) return "H"  ;
    if (arc_index == 1274) return "H"  ;
    if (arc_index == 1275) return "H"  ;
    if (arc_index == 1283) return "E"  ;
    if (arc_index == 1291) return "E"  ;
    if (arc_index == 1302) return "W"  ;
    if (arc_index == 1332) return "W"  ;
    if (arc_index == 1361) return "W"  ;
    if (arc_index == 1363) return "W"  ;
    if (arc_index == 1370) return "H"  ;
    if (arc_index == 1380) return "E"  ;
    if (arc_index == 1382) return "E"  ;
    if (arc_index == 1434) return "E"  ;
    if (arc_index == 1436) return "E"  ;
    if (arc_index == 1446) return "E"  ;
    if (arc_index == 1450) return "E"  ;
    if (arc_index == 1474) return "W"  ;
    if (arc_index == 1489) return "W"  ;
    if (arc_index == 1501) return "W"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1546) return "W"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1553) return "W"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1595) return "W"  ;
    if (arc_index == 1668) return "W"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1677) return "E"  ;
    if (arc_index == 1678) return "E"  ;
    if (arc_index == 1686) return "E"  ;
    if (arc_index == 1692) return "E"  ;
    if (arc_index == 1693) return "E"  ;
    if (arc_index == 1708) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1763) return "E"  ;
    if (arc_index == 1792) return "E"  ;
    if (arc_index == 1805) return "E"  ;
    if (arc_index == 1809) return "E"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1867) return "E"  ;
    if (arc_index == 1870) return "E"  ;
    if (arc_index == 1874) return "E"  ;
    if (arc_index == 1875) return "E"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1880) return "E"  ;
    if (arc_index == 1882) return "E"  ;
    if (arc_index == 1888) return "E"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1891) return "E"  ;
    if (arc_index == 1901) return "E"  ;
    if (arc_index == 1903) return "E"  ;
    if (arc_index == 1916) return "E"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1962) return "E"  ;
    if (arc_index == 1974) return "E"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2019) return "H"  ;
    if (arc_index == 2046) return "E"  ;
    if (arc_index == 2048) return "E"  ;
    if (arc_index == 2079) return "E"  ;
    if (arc_index == 2098) return "E"  ;
    if (arc_index == 2106) return "E"  ;
    if (arc_index == 2113) return "E"  ;
    if (arc_index == 2136) return "E"  ;
    if (arc_index == 2141) return "E"  ;
    if (arc_index == 2156) return "E"  ;
    if (arc_index == 2174) return "H"  ;
    if (arc_index == 2179) return "W"  ;
    if (arc_index == 2183) return "W"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2188) return "W"  ;
    if (arc_index == 2189) return "W"  ;
    if (arc_index == 2190) return "W"  ;
    if (arc_index == 2193) return "W"  ;
    if (arc_index == 2210) return "W"  ;
    if (arc_index == 2214) return "W"  ;
    if (arc_index == 2215) return "W"  ;
    if (arc_index == 2218) return "W"  ;
    if (arc_index == 2245) return "E"  ;
    if (arc_index == 2256) return "E"  ;
    if (arc_index == 2267) return "E"  ;
    if (arc_index == 2269) return "E"  ;
    if (arc_index == 2271) return "E"  ;
    if (arc_index == 2272) return "E"  ;
    if (arc_index == 2278) return "E"  ;
    if (arc_index == 2288) return "E"  ;
    if (arc_index == 2307) return "H"  ;
    if (arc_index == 2315) return "H"  ;
    if (arc_index == 2319) return "H"  ;
    if (arc_index == 2323) return "W"  ;
    if (arc_index == 2344) return "W"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2361) return "W"  ;
    if (arc_index == 2402) return "H"  ;
    if (arc_index == 2404) return "H"  ;
    if (arc_index == 2408) return "H"  ;
    if (arc_index == 2417) return "W"  ;
    if (arc_index == 2418) return "W"  ;
    if (arc_index == 2431) return "E"  ;
    if (arc_index == 2435) return "E"  ;
    if (arc_index == 2462) return "E"  ;
    if (arc_index == 2524) return "E"  ;
    if (arc_index == 2528) return "H"  ;
    if (arc_index == 2599) return "H"  ;
    if (arc_index == 2600) return "H"  ;
    if (arc_index == 2633) return "H"  ;
    if (arc_index == 2638) return "W"  ;
    if (arc_index == 2639) return "H"  ;
    if (arc_index == 2644) return "H"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2708) return "W"  ;
    if (arc_index == 2709) return "H"  ;
    if (arc_index == 2720) return "W"  ;
    if (arc_index == 2721) return "W"  ;
    if (arc_index == 2722) return "W"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2738) return "W"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2821) return "E"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2884) return "H"  ;
    if (arc_index == 2905) return "W"  ;
    if (arc_index == 2907) return "W"  ;
    if (arc_index == 2908) return "W"  ;
    if (arc_index == 2913) return "W"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 8)) begin 
    if (arc_index == 16) return "W"  ;
    if (arc_index == 30) return "W"  ;
    if (arc_index == 86) return "E"  ;
    if (arc_index == 161) return "E"  ;
    if (arc_index == 164) return "W"  ;
    if (arc_index == 177) return "H"  ;
    if (arc_index == 208) return "E"  ;
    if (arc_index == 220) return "H"  ;
    if (arc_index == 242) return "H"  ;
    if (arc_index == 243) return "E"  ;
    if (arc_index == 244) return "E"  ;
    if (arc_index == 245) return "E"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 247) return "W"  ;
    if (arc_index == 248) return "W"  ;
    if (arc_index == 249) return "W"  ;
    if (arc_index == 250) return "W"  ;
    if (arc_index == 251) return "W"  ;
    if (arc_index == 252) return "W"  ;
    if (arc_index == 253) return "W"  ;
    if (arc_index == 254) return "E"  ;
    if (arc_index == 255) return "E"  ;
    if (arc_index == 256) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 258) return "E"  ;
    if (arc_index == 259) return "W"  ;
    if (arc_index == 260) return "W"  ;
    if (arc_index == 261) return "W"  ;
    if (arc_index == 262) return "W"  ;
    if (arc_index == 263) return "W"  ;
    if (arc_index == 275) return "H"  ;
    if (arc_index == 320) return "H"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 519) return "H"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 528) return "E"  ;
    if (arc_index == 552) return "E"  ;
    if (arc_index == 556) return "E"  ;
    if (arc_index == 566) return "E"  ;
    if (arc_index == 568) return "E"  ;
    if (arc_index == 621) return "W"  ;
    if (arc_index == 683) return "W"  ;
    if (arc_index == 696) return "H"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 708) return "W"  ;
    if (arc_index == 710) return "W"  ;
    if (arc_index == 712) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 719) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 721) return "W"  ;
    if (arc_index == 722) return "W"  ;
    if (arc_index == 780) return "H"  ;
    if (arc_index == 782) return "E"  ;
    if (arc_index == 834) return "W"  ;
    if (arc_index == 889) return "H"  ;
    if (arc_index == 921) return "H"  ;
    if (arc_index == 929) return "H"  ;
    if (arc_index == 1005) return "H"  ;
    if (arc_index == 1016) return "H"  ;
    if (arc_index == 1094) return "H"  ;
    if (arc_index == 1108) return "H"  ;
    if (arc_index == 1118) return "H"  ;
    if (arc_index == 1146) return "W"  ;
    if (arc_index == 1239) return "H"  ;
    if (arc_index == 1251) return "H"  ;
    if (arc_index == 1259) return "H"  ;
    if (arc_index == 1392) return "H"  ;
    if (arc_index == 1420) return "H"  ;
    if (arc_index == 1426) return "H"  ;
    if (arc_index == 1458) return "H"  ;
    if (arc_index == 1467) return "E"  ;
    if (arc_index == 1468) return "E"  ;
    if (arc_index == 1469) return "E"  ;
    if (arc_index == 1583) return "E"  ;
    if (arc_index == 1624) return "E"  ;
    if (arc_index == 1653) return "E"  ;
    if (arc_index == 1685) return "W"  ;
    if (arc_index == 1701) return "E"  ;
    if (arc_index == 1705) return "E"  ;
    if (arc_index == 1708) return "E"  ;
    if (arc_index == 1738) return "E"  ;
    if (arc_index == 1757) return "E"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1760) return "W"  ;
    if (arc_index == 1763) return "W"  ;
    if (arc_index == 1764) return "W"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1773) return "W"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1778) return "W"  ;
    if (arc_index == 1781) return "W"  ;
    if (arc_index == 1793) return "W"  ;
    if (arc_index == 1828) return "W"  ;
    if (arc_index == 1854) return "E"  ;
    if (arc_index == 1978) return "E"  ;
    if (arc_index == 2041) return "H"  ;
    if (arc_index == 2068) return "H"  ;
    if (arc_index == 2090) return "H"  ;
    if (arc_index == 2091) return "H"  ;
    if (arc_index == 2092) return "E"  ;
    if (arc_index == 2093) return "E"  ;
    if (arc_index == 2095) return "E"  ;
    if (arc_index == 2097) return "E"  ;
    if (arc_index == 2098) return "E"  ;
    if (arc_index == 2100) return "E"  ;
    if (arc_index == 2103) return "E"  ;
    if (arc_index == 2104) return "E"  ;
    if (arc_index == 2106) return "E"  ;
    if (arc_index == 2108) return "E"  ;
    if (arc_index == 2123) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2196) return "H"  ;
    if (arc_index == 2214) return "H"  ;
    if (arc_index == 2289) return "E"  ;
    if (arc_index == 2329) return "H"  ;
    if (arc_index == 2337) return "H"  ;
    if (arc_index == 2341) return "W"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2367) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2424) return "H"  ;
    if (arc_index == 2503) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2531) return "E"  ;
    if (arc_index == 2550) return "H"  ;
    if (arc_index == 2572) return "H"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2602) return "W"  ;
    if (arc_index == 2603) return "W"  ;
    if (arc_index == 2604) return "W"  ;
    if (arc_index == 2605) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2608) return "W"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2617) return "W"  ;
    if (arc_index == 2661) return "H"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2731) return "H"  ;
    if (arc_index == 2791) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2873) return "E"  ;
    if (arc_index == 2906) return "H"  ;
    if (arc_index == 2916) return "H"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 8)) begin 
    if (arc_index == 2) return "H"  ;
    if (arc_index == 8) return "E"  ;
    if (arc_index == 10) return "E"  ;
    if (arc_index == 11) return "E"  ;
    if (arc_index == 15) return "E"  ;
    if (arc_index == 17) return "E"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 89) return "E"  ;
    if (arc_index == 97) return "E"  ;
    if (arc_index == 109) return "E"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 154) return "E"  ;
    if (arc_index == 155) return "E"  ;
    if (arc_index == 156) return "W"  ;
    if (arc_index == 157) return "E"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 163) return "W"  ;
    if (arc_index == 165) return "W"  ;
    if (arc_index == 166) return "W"  ;
    if (arc_index == 170) return "W"  ;
    if (arc_index == 171) return "W"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 177) return "W"  ;
    if (arc_index == 187) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 198) return "W"  ;
    if (arc_index == 199) return "H"  ;
    if (arc_index == 209) return "H"  ;
    if (arc_index == 219) return "H"  ;
    if (arc_index == 220) return "H"  ;
    if (arc_index == 225) return "W"  ;
    if (arc_index == 228) return "W"  ;
    if (arc_index == 231) return "W"  ;
    if (arc_index == 232) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 242) return "H"  ;
    if (arc_index == 249) return "H"  ;
    if (arc_index == 250) return "H"  ;
    if (arc_index == 252) return "H"  ;
    if (arc_index == 253) return "H"  ;
    if (arc_index == 260) return "H"  ;
    if (arc_index == 264) return "E"  ;
    if (arc_index == 265) return "W"  ;
    if (arc_index == 266) return "E"  ;
    if (arc_index == 267) return "E"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 269) return "W"  ;
    if (arc_index == 270) return "W"  ;
    if (arc_index == 271) return "W"  ;
    if (arc_index == 272) return "E"  ;
    if (arc_index == 273) return "E"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 275) return "W"  ;
    if (arc_index == 276) return "W"  ;
    if (arc_index == 277) return "W"  ;
    if (arc_index == 278) return "W"  ;
    if (arc_index == 279) return "W"  ;
    if (arc_index == 280) return "E"  ;
    if (arc_index == 281) return "E"  ;
    if (arc_index == 282) return "E"  ;
    if (arc_index == 283) return "E"  ;
    if (arc_index == 284) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 296) return "W"  ;
    if (arc_index == 297) return "H"  ;
    if (arc_index == 321) return "H"  ;
    if (arc_index == 332) return "E"  ;
    if (arc_index == 342) return "H"  ;
    if (arc_index == 400) return "H"  ;
    if (arc_index == 420) return "H"  ;
    if (arc_index == 431) return "H"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 481) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 538) return "W"  ;
    if (arc_index == 541) return "H"  ;
    if (arc_index == 547) return "H"  ;
    if (arc_index == 549) return "W"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 595) return "W"  ;
    if (arc_index == 599) return "W"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 603) return "W"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 607) return "W"  ;
    if (arc_index == 609) return "W"  ;
    if (arc_index == 610) return "W"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 619) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 643) return "W"  ;
    if (arc_index == 660) return "W"  ;
    if (arc_index == 667) return "W"  ;
    if (arc_index == 695) return "W"  ;
    if (arc_index == 700) return "W"  ;
    if (arc_index == 702) return "E"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 718) return "H"  ;
    if (arc_index == 730) return "H"  ;
    if (arc_index == 758) return "H"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 802) return "H"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 833) return "W"  ;
    if (arc_index == 841) return "W"  ;
    if (arc_index == 883) return "E"  ;
    if (arc_index == 911) return "H"  ;
    if (arc_index == 917) return "H"  ;
    if (arc_index == 929) return "H"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1027) return "H"  ;
    if (arc_index == 1034) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1040) return "W"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1058) return "E"  ;
    if (arc_index == 1066) return "E"  ;
    if (arc_index == 1067) return "E"  ;
    if (arc_index == 1071) return "E"  ;
    if (arc_index == 1116) return "H"  ;
    if (arc_index == 1130) return "H"  ;
    if (arc_index == 1133) return "W"  ;
    if (arc_index == 1134) return "W"  ;
    if (arc_index == 1136) return "W"  ;
    if (arc_index == 1144) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1148) return "W"  ;
    if (arc_index == 1150) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1165) return "W"  ;
    if (arc_index == 1177) return "W"  ;
    if (arc_index == 1222) return "W"  ;
    if (arc_index == 1227) return "W"  ;
    if (arc_index == 1236) return "W"  ;
    if (arc_index == 1239) return "W"  ;
    if (arc_index == 1251) return "W"  ;
    if (arc_index == 1257) return "W"  ;
    if (arc_index == 1259) return "W"  ;
    if (arc_index == 1261) return "H"  ;
    if (arc_index == 1263) return "H"  ;
    if (arc_index == 1304) return "H"  ;
    if (arc_index == 1321) return "W"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1325) return "W"  ;
    if (arc_index == 1327) return "W"  ;
    if (arc_index == 1328) return "W"  ;
    if (arc_index == 1329) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1332) return "W"  ;
    if (arc_index == 1333) return "W"  ;
    if (arc_index == 1334) return "W"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1341) return "W"  ;
    if (arc_index == 1354) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1363) return "W"  ;
    if (arc_index == 1375) return "E"  ;
    if (arc_index == 1398) return "E"  ;
    if (arc_index == 1410) return "E"  ;
    if (arc_index == 1414) return "H"  ;
    if (arc_index == 1445) return "H"  ;
    if (arc_index == 1460) return "E"  ;
    if (arc_index == 1474) return "E"  ;
    if (arc_index == 1479) return "E"  ;
    if (arc_index == 1480) return "W"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1488) return "W"  ;
    if (arc_index == 1489) return "W"  ;
    if (arc_index == 1490) return "W"  ;
    if (arc_index == 1501) return "W"  ;
    if (arc_index == 1507) return "W"  ;
    if (arc_index == 1523) return "W"  ;
    if (arc_index == 1544) return "W"  ;
    if (arc_index == 1554) return "W"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1672) return "W"  ;
    if (arc_index == 1673) return "W"  ;
    if (arc_index == 1679) return "W"  ;
    if (arc_index == 1680) return "W"  ;
    if (arc_index == 1682) return "E"  ;
    if (arc_index == 1685) return "E"  ;
    if (arc_index == 1688) return "E"  ;
    if (arc_index == 1689) return "W"  ;
    if (arc_index == 1705) return "W"  ;
    if (arc_index == 1708) return "W"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1763) return "E"  ;
    if (arc_index == 1792) return "E"  ;
    if (arc_index == 1805) return "E"  ;
    if (arc_index == 1806) return "E"  ;
    if (arc_index == 1809) return "E"  ;
    if (arc_index == 1858) return "E"  ;
    if (arc_index == 1867) return "E"  ;
    if (arc_index == 1882) return "E"  ;
    if (arc_index == 1888) return "E"  ;
    if (arc_index == 1903) return "E"  ;
    if (arc_index == 1907) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1953) return "E"  ;
    if (arc_index == 1964) return "E"  ;
    if (arc_index == 1967) return "E"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 2063) return "H"  ;
    if (arc_index == 2072) return "H"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2081) return "W"  ;
    if (arc_index == 2098) return "W"  ;
    if (arc_index == 2106) return "W"  ;
    if (arc_index == 2182) return "W"  ;
    if (arc_index == 2214) return "W"  ;
    if (arc_index == 2215) return "W"  ;
    if (arc_index == 2218) return "H"  ;
    if (arc_index == 2249) return "H"  ;
    if (arc_index == 2267) return "E"  ;
    if (arc_index == 2286) return "E"  ;
    if (arc_index == 2307) return "E"  ;
    if (arc_index == 2313) return "E"  ;
    if (arc_index == 2320) return "W"  ;
    if (arc_index == 2329) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2344) return "W"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2351) return "H"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2359) return "H"  ;
    if (arc_index == 2372) return "H"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2386) return "W"  ;
    if (arc_index == 2389) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2413) return "W"  ;
    if (arc_index == 2419) return "W"  ;
    if (arc_index == 2446) return "H"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2462) return "E"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2470) return "E"  ;
    if (arc_index == 2476) return "E"  ;
    if (arc_index == 2482) return "E"  ;
    if (arc_index == 2537) return "E"  ;
    if (arc_index == 2538) return "E"  ;
    if (arc_index == 2548) return "E"  ;
    if (arc_index == 2572) return "H"  ;
    if (arc_index == 2599) return "H"  ;
    if (arc_index == 2600) return "H"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2683) return "H"  ;
    if (arc_index == 2689) return "E"  ;
    if (arc_index == 2690) return "E"  ;
    if (arc_index == 2696) return "E"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2753) return "H"  ;
    if (arc_index == 2784) return "H"  ;
    if (arc_index == 2822) return "H"  ;
    if (arc_index == 2825) return "E"  ;
    if (arc_index == 2831) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2895) return "E"  ;
    if (arc_index == 2902) return "E"  ;
    if (arc_index == 2904) return "W"  ;
    if (arc_index == 2907) return "W"  ;
    if (arc_index == 2913) return "W"  ;
    if (arc_index == 2922) return "W"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 10)) begin 
    if (arc_index == 15) return "W"  ;
    if (arc_index == 24) return "H"  ;
    if (arc_index == 168) return "E"  ;
    if (arc_index == 179) return "E"  ;
    if (arc_index == 191) return "E"  ;
    if (arc_index == 196) return "W"  ;
    if (arc_index == 197) return "W"  ;
    if (arc_index == 203) return "W"  ;
    if (arc_index == 221) return "H"  ;
    if (arc_index == 230) return "E"  ;
    if (arc_index == 254) return "E"  ;
    if (arc_index == 264) return "H"  ;
    if (arc_index == 286) return "H"  ;
    if (arc_index == 287) return "H"  ;
    if (arc_index == 288) return "H"  ;
    if (arc_index == 289) return "H"  ;
    if (arc_index == 290) return "H"  ;
    if (arc_index == 291) return "H"  ;
    if (arc_index == 292) return "H"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 294) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 296) return "W"  ;
    if (arc_index == 297) return "W"  ;
    if (arc_index == 298) return "W"  ;
    if (arc_index == 299) return "W"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 301) return "W"  ;
    if (arc_index == 302) return "W"  ;
    if (arc_index == 303) return "W"  ;
    if (arc_index == 304) return "W"  ;
    if (arc_index == 305) return "W"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 307) return "W"  ;
    if (arc_index == 319) return "H"  ;
    if (arc_index == 364) return "H"  ;
    if (arc_index == 370) return "H"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 544) return "E"  ;
    if (arc_index == 563) return "H"  ;
    if (arc_index == 566) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 597) return "E"  ;
    if (arc_index == 614) return "E"  ;
    if (arc_index == 615) return "E"  ;
    if (arc_index == 616) return "E"  ;
    if (arc_index == 620) return "E"  ;
    if (arc_index == 630) return "E"  ;
    if (arc_index == 636) return "W"  ;
    if (arc_index == 639) return "W"  ;
    if (arc_index == 672) return "W"  ;
    if (arc_index == 701) return "E"  ;
    if (arc_index == 714) return "E"  ;
    if (arc_index == 723) return "E"  ;
    if (arc_index == 740) return "H"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 824) return "H"  ;
    if (arc_index == 871) return "H"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 933) return "H"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1034) return "E"  ;
    if (arc_index == 1037) return "W"  ;
    if (arc_index == 1048) return "W"  ;
    if (arc_index == 1049) return "H"  ;
    if (arc_index == 1054) return "W"  ;
    if (arc_index == 1067) return "W"  ;
    if (arc_index == 1122) return "W"  ;
    if (arc_index == 1128) return "E"  ;
    if (arc_index == 1132) return "E"  ;
    if (arc_index == 1138) return "H"  ;
    if (arc_index == 1141) return "H"  ;
    if (arc_index == 1152) return "H"  ;
    if (arc_index == 1155) return "H"  ;
    if (arc_index == 1163) return "H"  ;
    if (arc_index == 1241) return "H"  ;
    if (arc_index == 1242) return "H"  ;
    if (arc_index == 1249) return "E"  ;
    if (arc_index == 1277) return "E"  ;
    if (arc_index == 1278) return "E"  ;
    if (arc_index == 1283) return "H"  ;
    if (arc_index == 1305) return "H"  ;
    if (arc_index == 1326) return "H"  ;
    if (arc_index == 1339) return "H"  ;
    if (arc_index == 1342) return "H"  ;
    if (arc_index == 1347) return "H"  ;
    if (arc_index == 1361) return "W"  ;
    if (arc_index == 1436) return "H"  ;
    if (arc_index == 1446) return "H"  ;
    if (arc_index == 1475) return "E"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1541) return "W"  ;
    if (arc_index == 1542) return "W"  ;
    if (arc_index == 1543) return "W"  ;
    if (arc_index == 1544) return "W"  ;
    if (arc_index == 1546) return "W"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1553) return "W"  ;
    if (arc_index == 1554) return "W"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1559) return "W"  ;
    if (arc_index == 1560) return "W"  ;
    if (arc_index == 1570) return "W"  ;
    if (arc_index == 1577) return "W"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1681) return "E"  ;
    if (arc_index == 1769) return "E"  ;
    if (arc_index == 1806) return "E"  ;
    if (arc_index == 1874) return "E"  ;
    if (arc_index == 1994) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2075) return "E"  ;
    if (arc_index == 2081) return "E"  ;
    if (arc_index == 2083) return "W"  ;
    if (arc_index == 2085) return "H"  ;
    if (arc_index == 2089) return "H"  ;
    if (arc_index == 2101) return "H"  ;
    if (arc_index == 2114) return "E"  ;
    if (arc_index == 2181) return "E"  ;
    if (arc_index == 2182) return "W"  ;
    if (arc_index == 2187) return "E"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2194) return "W"  ;
    if (arc_index == 2196) return "W"  ;
    if (arc_index == 2198) return "W"  ;
    if (arc_index == 2208) return "W"  ;
    if (arc_index == 2240) return "H"  ;
    if (arc_index == 2303) return "E"  ;
    if (arc_index == 2311) return "E"  ;
    if (arc_index == 2345) return "E"  ;
    if (arc_index == 2358) return "E"  ;
    if (arc_index == 2373) return "H"  ;
    if (arc_index == 2376) return "W"  ;
    if (arc_index == 2377) return "W"  ;
    if (arc_index == 2381) return "H"  ;
    if (arc_index == 2382) return "H"  ;
    if (arc_index == 2406) return "E"  ;
    if (arc_index == 2409) return "E"  ;
    if (arc_index == 2468) return "H"  ;
    if (arc_index == 2484) return "H"  ;
    if (arc_index == 2537) return "E"  ;
    if (arc_index == 2594) return "H"  ;
    if (arc_index == 2606) return "H"  ;
    if (arc_index == 2623) return "W"  ;
    if (arc_index == 2632) return "W"  ;
    if (arc_index == 2633) return "W"  ;
    if (arc_index == 2638) return "W"  ;
    if (arc_index == 2639) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2690) return "E"  ;
    if (arc_index == 2705) return "H"  ;
    if (arc_index == 2775) return "H"  ;
    if (arc_index == 2825) return "H"  ;
    if (arc_index == 2833) return "E"  ;
    if (arc_index == 2905) return "W"  ;
    if (arc_index == 2908) return "W"  ;
    if (arc_index == 2920) return "W"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 10)) begin 
    if (arc_index == 46) return "H"  ;
    if (arc_index == 109) return "E"  ;
    if (arc_index == 197) return "E"  ;
    if (arc_index == 243) return "H"  ;
    if (arc_index == 254) return "H"  ;
    if (arc_index == 267) return "H"  ;
    if (arc_index == 286) return "H"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 308) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 311) return "W"  ;
    if (arc_index == 312) return "W"  ;
    if (arc_index == 313) return "W"  ;
    if (arc_index == 314) return "W"  ;
    if (arc_index == 315) return "W"  ;
    if (arc_index == 316) return "W"  ;
    if (arc_index == 317) return "W"  ;
    if (arc_index == 318) return "W"  ;
    if (arc_index == 319) return "W"  ;
    if (arc_index == 320) return "W"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 323) return "W"  ;
    if (arc_index == 324) return "W"  ;
    if (arc_index == 325) return "W"  ;
    if (arc_index == 326) return "W"  ;
    if (arc_index == 327) return "W"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 329) return "W"  ;
    if (arc_index == 341) return "H"  ;
    if (arc_index == 354) return "E"  ;
    if (arc_index == 386) return "H"  ;
    if (arc_index == 558) return "E"  ;
    if (arc_index == 563) return "E"  ;
    if (arc_index == 585) return "H"  ;
    if (arc_index == 617) return "W"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 619) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 627) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 634) return "W"  ;
    if (arc_index == 635) return "W"  ;
    if (arc_index == 639) return "W"  ;
    if (arc_index == 649) return "E"  ;
    if (arc_index == 694) return "E"  ;
    if (arc_index == 704) return "E"  ;
    if (arc_index == 706) return "E"  ;
    if (arc_index == 707) return "E"  ;
    if (arc_index == 709) return "E"  ;
    if (arc_index == 711) return "E"  ;
    if (arc_index == 714) return "E"  ;
    if (arc_index == 716) return "E"  ;
    if (arc_index == 718) return "E"  ;
    if (arc_index == 723) return "E"  ;
    if (arc_index == 724) return "E"  ;
    if (arc_index == 725) return "E"  ;
    if (arc_index == 737) return "E"  ;
    if (arc_index == 762) return "H"  ;
    if (arc_index == 846) return "H"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 955) return "H"  ;
    if (arc_index == 981) return "H"  ;
    if (arc_index == 1070) return "E"  ;
    if (arc_index == 1071) return "H"  ;
    if (arc_index == 1158) return "H"  ;
    if (arc_index == 1160) return "H"  ;
    if (arc_index == 1174) return "H"  ;
    if (arc_index == 1242) return "H"  ;
    if (arc_index == 1263) return "E"  ;
    if (arc_index == 1305) return "H"  ;
    if (arc_index == 1346) return "H"  ;
    if (arc_index == 1351) return "H"  ;
    if (arc_index == 1360) return "W"  ;
    if (arc_index == 1379) return "E"  ;
    if (arc_index == 1458) return "H"  ;
    if (arc_index == 1468) return "E"  ;
    if (arc_index == 1547) return "E"  ;
    if (arc_index == 1548) return "W"  ;
    if (arc_index == 1556) return "W"  ;
    if (arc_index == 1570) return "W"  ;
    if (arc_index == 1613) return "E"  ;
    if (arc_index == 1766) return "E"  ;
    if (arc_index == 2101) return "E"  ;
    if (arc_index == 2105) return "E"  ;
    if (arc_index == 2107) return "H"  ;
    if (arc_index == 2111) return "E"  ;
    if (arc_index == 2262) return "H"  ;
    if (arc_index == 2339) return "H"  ;
    if (arc_index == 2380) return "W"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2395) return "H"  ;
    if (arc_index == 2403) return "H"  ;
    if (arc_index == 2490) return "H"  ;
    if (arc_index == 2553) return "H"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2596) return "E"  ;
    if (arc_index == 2616) return "H"  ;
    if (arc_index == 2626) return "H"  ;
    if (arc_index == 2628) return "H"  ;
    if (arc_index == 2629) return "H"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2635) return "W"  ;
    if (arc_index == 2636) return "W"  ;
    if (arc_index == 2637) return "W"  ;
    if (arc_index == 2658) return "W"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2727) return "H"  ;
    if (arc_index == 2797) return "H"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2906) return "W"  ;
    if (arc_index == 2916) return "W"  ;
    if (arc_index == 2923) return "W"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 6)) begin 
    if (arc_index == 1) return "W"  ;
    if (arc_index == 3) return "W"  ;
    if (arc_index == 19) return "W"  ;
    if (arc_index == 20) return "W"  ;
    if (arc_index == 29) return "E"  ;
    if (arc_index == 33) return "E"  ;
    if (arc_index == 43) return "E"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 53) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 57) return "E"  ;
    if (arc_index == 62) return "E"  ;
    if (arc_index == 68) return "H"  ;
    if (arc_index == 98) return "H"  ;
    if (arc_index == 113) return "H"  ;
    if (arc_index == 119) return "E"  ;
    if (arc_index == 128) return "E"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 165) return "E"  ;
    if (arc_index == 173) return "E"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 184) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 201) return "W"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 222) return "W"  ;
    if (arc_index == 223) return "W"  ;
    if (arc_index == 224) return "W"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 227) return "W"  ;
    if (arc_index == 238) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 265) return "H"  ;
    if (arc_index == 299) return "H"  ;
    if (arc_index == 303) return "W"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 308) return "H"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 327) return "W"  ;
    if (arc_index == 330) return "W"  ;
    if (arc_index == 331) return "W"  ;
    if (arc_index == 332) return "W"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 335) return "W"  ;
    if (arc_index == 336) return "W"  ;
    if (arc_index == 337) return "E"  ;
    if (arc_index == 338) return "E"  ;
    if (arc_index == 339) return "E"  ;
    if (arc_index == 340) return "E"  ;
    if (arc_index == 341) return "E"  ;
    if (arc_index == 342) return "E"  ;
    if (arc_index == 343) return "W"  ;
    if (arc_index == 344) return "W"  ;
    if (arc_index == 345) return "W"  ;
    if (arc_index == 346) return "W"  ;
    if (arc_index == 347) return "W"  ;
    if (arc_index == 348) return "E"  ;
    if (arc_index == 349) return "W"  ;
    if (arc_index == 350) return "W"  ;
    if (arc_index == 351) return "W"  ;
    if (arc_index == 356) return "W"  ;
    if (arc_index == 363) return "H"  ;
    if (arc_index == 373) return "H"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 402) return "E"  ;
    if (arc_index == 408) return "H"  ;
    if (arc_index == 426) return "H"  ;
    if (arc_index == 436) return "H"  ;
    if (arc_index == 490) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 497) return "E"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 530) return "W"  ;
    if (arc_index == 540) return "W"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 564) return "W"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 599) return "W"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 607) return "H"  ;
    if (arc_index == 629) return "H"  ;
    if (arc_index == 639) return "E"  ;
    if (arc_index == 642) return "E"  ;
    if (arc_index == 647) return "E"  ;
    if (arc_index == 649) return "E"  ;
    if (arc_index == 653) return "E"  ;
    if (arc_index == 654) return "E"  ;
    if (arc_index == 655) return "E"  ;
    if (arc_index == 656) return "E"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 674) return "E"  ;
    if (arc_index == 677) return "E"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 769) return "E"  ;
    if (arc_index == 784) return "H"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 836) return "E"  ;
    if (arc_index == 839) return "E"  ;
    if (arc_index == 850) return "E"  ;
    if (arc_index == 851) return "E"  ;
    if (arc_index == 863) return "E"  ;
    if (arc_index == 866) return "E"  ;
    if (arc_index == 868) return "H"  ;
    if (arc_index == 869) return "H"  ;
    if (arc_index == 876) return "H"  ;
    if (arc_index == 890) return "H"  ;
    if (arc_index == 898) return "H"  ;
    if (arc_index == 904) return "H"  ;
    if (arc_index == 928) return "H"  ;
    if (arc_index == 929) return "H"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 973) return "E"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 977) return "H"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 983) return "E"  ;
    if (arc_index == 986) return "E"  ;
    if (arc_index == 997) return "E"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1044) return "E"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1059) return "W"  ;
    if (arc_index == 1085) return "W"  ;
    if (arc_index == 1092) return "W"  ;
    if (arc_index == 1093) return "H"  ;
    if (arc_index == 1100) return "H"  ;
    if (arc_index == 1101) return "H"  ;
    if (arc_index == 1102) return "H"  ;
    if (arc_index == 1107) return "H"  ;
    if (arc_index == 1114) return "H"  ;
    if (arc_index == 1115) return "H"  ;
    if (arc_index == 1143) return "H"  ;
    if (arc_index == 1168) return "W"  ;
    if (arc_index == 1170) return "W"  ;
    if (arc_index == 1174) return "W"  ;
    if (arc_index == 1175) return "E"  ;
    if (arc_index == 1177) return "E"  ;
    if (arc_index == 1178) return "E"  ;
    if (arc_index == 1182) return "H"  ;
    if (arc_index == 1185) return "H"  ;
    if (arc_index == 1186) return "H"  ;
    if (arc_index == 1187) return "H"  ;
    if (arc_index == 1196) return "H"  ;
    if (arc_index == 1212) return "H"  ;
    if (arc_index == 1214) return "E"  ;
    if (arc_index == 1217) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1250) return "E"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1272) return "W"  ;
    if (arc_index == 1279) return "W"  ;
    if (arc_index == 1281) return "W"  ;
    if (arc_index == 1292) return "W"  ;
    if (arc_index == 1296) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1325) return "W"  ;
    if (arc_index == 1327) return "H"  ;
    if (arc_index == 1349) return "H"  ;
    if (arc_index == 1368) return "W"  ;
    if (arc_index == 1377) return "W"  ;
    if (arc_index == 1385) return "W"  ;
    if (arc_index == 1396) return "W"  ;
    if (arc_index == 1397) return "E"  ;
    if (arc_index == 1401) return "E"  ;
    if (arc_index == 1415) return "E"  ;
    if (arc_index == 1434) return "E"  ;
    if (arc_index == 1435) return "E"  ;
    if (arc_index == 1436) return "E"  ;
    if (arc_index == 1443) return "E"  ;
    if (arc_index == 1445) return "E"  ;
    if (arc_index == 1446) return "E"  ;
    if (arc_index == 1449) return "E"  ;
    if (arc_index == 1450) return "E"  ;
    if (arc_index == 1451) return "E"  ;
    if (arc_index == 1456) return "E"  ;
    if (arc_index == 1462) return "W"  ;
    if (arc_index == 1471) return "W"  ;
    if (arc_index == 1474) return "W"  ;
    if (arc_index == 1480) return "H"  ;
    if (arc_index == 1490) return "H"  ;
    if (arc_index == 1500) return "H"  ;
    if (arc_index == 1507) return "H"  ;
    if (arc_index == 1515) return "E"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1522) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1551) return "E"  ;
    if (arc_index == 1608) return "E"  ;
    if (arc_index == 1620) return "E"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1641) return "E"  ;
    if (arc_index == 1648) return "E"  ;
    if (arc_index == 1687) return "E"  ;
    if (arc_index == 1704) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1764) return "E"  ;
    if (arc_index == 1788) return "E"  ;
    if (arc_index == 1813) return "E"  ;
    if (arc_index == 1820) return "E"  ;
    if (arc_index == 1821) return "W"  ;
    if (arc_index == 1848) return "E"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1896) return "W"  ;
    if (arc_index == 1900) return "E"  ;
    if (arc_index == 1916) return "E"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1965) return "E"  ;
    if (arc_index == 1968) return "W"  ;
    if (arc_index == 1988) return "W"  ;
    if (arc_index == 2004) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2032) return "E"  ;
    if (arc_index == 2048) return "E"  ;
    if (arc_index == 2077) return "W"  ;
    if (arc_index == 2113) return "E"  ;
    if (arc_index == 2120) return "E"  ;
    if (arc_index == 2127) return "E"  ;
    if (arc_index == 2128) return "E"  ;
    if (arc_index == 2129) return "H"  ;
    if (arc_index == 2133) return "H"  ;
    if (arc_index == 2156) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2174) return "E"  ;
    if (arc_index == 2179) return "E"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2189) return "W"  ;
    if (arc_index == 2190) return "W"  ;
    if (arc_index == 2193) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2233) return "W"  ;
    if (arc_index == 2245) return "E"  ;
    if (arc_index == 2246) return "E"  ;
    if (arc_index == 2251) return "E"  ;
    if (arc_index == 2256) return "E"  ;
    if (arc_index == 2259) return "W"  ;
    if (arc_index == 2263) return "E"  ;
    if (arc_index == 2274) return "E"  ;
    if (arc_index == 2275) return "W"  ;
    if (arc_index == 2276) return "W"  ;
    if (arc_index == 2277) return "W"  ;
    if (arc_index == 2279) return "W"  ;
    if (arc_index == 2280) return "W"  ;
    if (arc_index == 2281) return "W"  ;
    if (arc_index == 2282) return "W"  ;
    if (arc_index == 2283) return "W"  ;
    if (arc_index == 2284) return "H"  ;
    if (arc_index == 2296) return "W"  ;
    if (arc_index == 2306) return "W"  ;
    if (arc_index == 2398) return "W"  ;
    if (arc_index == 2417) return "H"  ;
    if (arc_index == 2425) return "H"  ;
    if (arc_index == 2431) return "E"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2505) return "E"  ;
    if (arc_index == 2512) return "H"  ;
    if (arc_index == 2521) return "H"  ;
    if (arc_index == 2534) return "H"  ;
    if (arc_index == 2614) return "H"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2638) return "H"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2708) return "W"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2736) return "W"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2749) return "H"  ;
    if (arc_index == 2752) return "H"  ;
    if (arc_index == 2764) return "E"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2819) return "H"  ;
    if (arc_index == 2820) return "H"  ;
    if (arc_index == 2841) return "H"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2884) return "E"  ;
    if (arc_index == 2905) return "W"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 6)) begin 
    if (arc_index == 19) return "W"  ;
    if (arc_index == 37) return "E"  ;
    if (arc_index == 90) return "H"  ;
    if (arc_index == 114) return "H"  ;
    if (arc_index == 140) return "E"  ;
    if (arc_index == 223) return "W"  ;
    if (arc_index == 287) return "H"  ;
    if (arc_index == 330) return "H"  ;
    if (arc_index == 351) return "H"  ;
    if (arc_index == 352) return "W"  ;
    if (arc_index == 353) return "E"  ;
    if (arc_index == 354) return "E"  ;
    if (arc_index == 355) return "W"  ;
    if (arc_index == 356) return "W"  ;
    if (arc_index == 357) return "W"  ;
    if (arc_index == 358) return "W"  ;
    if (arc_index == 359) return "W"  ;
    if (arc_index == 360) return "W"  ;
    if (arc_index == 361) return "E"  ;
    if (arc_index == 362) return "E"  ;
    if (arc_index == 363) return "E"  ;
    if (arc_index == 364) return "E"  ;
    if (arc_index == 365) return "E"  ;
    if (arc_index == 366) return "E"  ;
    if (arc_index == 367) return "E"  ;
    if (arc_index == 368) return "W"  ;
    if (arc_index == 369) return "W"  ;
    if (arc_index == 370) return "E"  ;
    if (arc_index == 371) return "E"  ;
    if (arc_index == 372) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 385) return "H"  ;
    if (arc_index == 392) return "H"  ;
    if (arc_index == 416) return "E"  ;
    if (arc_index == 418) return "W"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 429) return "W"  ;
    if (arc_index == 430) return "H"  ;
    if (arc_index == 434) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 595) return "E"  ;
    if (arc_index == 596) return "E"  ;
    if (arc_index == 629) return "H"  ;
    if (arc_index == 638) return "W"  ;
    if (arc_index == 657) return "W"  ;
    if (arc_index == 660) return "W"  ;
    if (arc_index == 671) return "W"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 806) return "H"  ;
    if (arc_index == 813) return "H"  ;
    if (arc_index == 825) return "W"  ;
    if (arc_index == 836) return "W"  ;
    if (arc_index == 862) return "W"  ;
    if (arc_index == 863) return "W"  ;
    if (arc_index == 866) return "W"  ;
    if (arc_index == 868) return "W"  ;
    if (arc_index == 869) return "W"  ;
    if (arc_index == 873) return "W"  ;
    if (arc_index == 874) return "W"  ;
    if (arc_index == 876) return "W"  ;
    if (arc_index == 879) return "W"  ;
    if (arc_index == 890) return "H"  ;
    if (arc_index == 891) return "H"  ;
    if (arc_index == 927) return "H"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 992) return "E"  ;
    if (arc_index == 999) return "H"  ;
    if (arc_index == 1003) return "E"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1041) return "W"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1069) return "W"  ;
    if (arc_index == 1114) return "W"  ;
    if (arc_index == 1115) return "H"  ;
    if (arc_index == 1123) return "W"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1171) return "W"  ;
    if (arc_index == 1180) return "E"  ;
    if (arc_index == 1181) return "E"  ;
    if (arc_index == 1204) return "H"  ;
    if (arc_index == 1218) return "H"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1234) return "W"  ;
    if (arc_index == 1246) return "W"  ;
    if (arc_index == 1312) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1315) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1349) return "H"  ;
    if (arc_index == 1365) return "H"  ;
    if (arc_index == 1368) return "H"  ;
    if (arc_index == 1383) return "H"  ;
    if (arc_index == 1396) return "H"  ;
    if (arc_index == 1456) return "E"  ;
    if (arc_index == 1497) return "E"  ;
    if (arc_index == 1501) return "E"  ;
    if (arc_index == 1502) return "H"  ;
    if (arc_index == 1505) return "H"  ;
    if (arc_index == 1510) return "E"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1574) return "W"  ;
    if (arc_index == 1621) return "W"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1723) return "E"  ;
    if (arc_index == 1810) return "W"  ;
    if (arc_index == 2017) return "E"  ;
    if (arc_index == 2018) return "E"  ;
    if (arc_index == 2019) return "E"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2119) return "E"  ;
    if (arc_index == 2135) return "E"  ;
    if (arc_index == 2150) return "E"  ;
    if (arc_index == 2151) return "H"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2180) return "W"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2204) return "W"  ;
    if (arc_index == 2212) return "W"  ;
    if (arc_index == 2219) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2306) return "H"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2377) return "W"  ;
    if (arc_index == 2439) return "H"  ;
    if (arc_index == 2444) return "E"  ;
    if (arc_index == 2447) return "H"  ;
    if (arc_index == 2448) return "E"  ;
    if (arc_index == 2455) return "E"  ;
    if (arc_index == 2462) return "E"  ;
    if (arc_index == 2513) return "E"  ;
    if (arc_index == 2534) return "H"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2577) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2614) return "E"  ;
    if (arc_index == 2646) return "W"  ;
    if (arc_index == 2660) return "H"  ;
    if (arc_index == 2673) return "H"  ;
    if (arc_index == 2771) return "H"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2841) return "H"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 1)) begin 
    if (arc_index == 112) return "H"  ;
    if (arc_index == 135) return "H"  ;
    if (arc_index == 268) return "H"  ;
    if (arc_index == 309) return "H"  ;
    if (arc_index == 352) return "H"  ;
    if (arc_index == 374) return "E"  ;
    if (arc_index == 375) return "E"  ;
    if (arc_index == 376) return "E"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 379) return "E"  ;
    if (arc_index == 380) return "E"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 382) return "E"  ;
    if (arc_index == 383) return "W"  ;
    if (arc_index == 384) return "W"  ;
    if (arc_index == 385) return "E"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 387) return "E"  ;
    if (arc_index == 388) return "E"  ;
    if (arc_index == 389) return "E"  ;
    if (arc_index == 390) return "E"  ;
    if (arc_index == 391) return "E"  ;
    if (arc_index == 392) return "E"  ;
    if (arc_index == 393) return "E"  ;
    if (arc_index == 394) return "E"  ;
    if (arc_index == 395) return "E"  ;
    if (arc_index == 407) return "H"  ;
    if (arc_index == 418) return "H"  ;
    if (arc_index == 452) return "H"  ;
    if (arc_index == 487) return "E"  ;
    if (arc_index == 505) return "E"  ;
    if (arc_index == 513) return "E"  ;
    if (arc_index == 514) return "E"  ;
    if (arc_index == 575) return "E"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 651) return "H"  ;
    if (arc_index == 750) return "H"  ;
    if (arc_index == 828) return "H"  ;
    if (arc_index == 912) return "H"  ;
    if (arc_index == 947) return "H"  ;
    if (arc_index == 1013) return "H"  ;
    if (arc_index == 1016) return "H"  ;
    if (arc_index == 1017) return "H"  ;
    if (arc_index == 1018) return "H"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1021) return "H"  ;
    if (arc_index == 1022) return "W"  ;
    if (arc_index == 1024) return "W"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1026) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1029) return "E"  ;
    if (arc_index == 1032) return "E"  ;
    if (arc_index == 1090) return "E"  ;
    if (arc_index == 1137) return "H"  ;
    if (arc_index == 1226) return "H"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1240) return "H"  ;
    if (arc_index == 1371) return "H"  ;
    if (arc_index == 1466) return "H"  ;
    if (arc_index == 1524) return "H"  ;
    if (arc_index == 1526) return "H"  ;
    if (arc_index == 1536) return "E"  ;
    if (arc_index == 1562) return "E"  ;
    if (arc_index == 1602) return "E"  ;
    if (arc_index == 1659) return "E"  ;
    if (arc_index == 1735) return "E"  ;
    if (arc_index == 1743) return "E"  ;
    if (arc_index == 1830) return "E"  ;
    if (arc_index == 1864) return "E"  ;
    if (arc_index == 1878) return "E"  ;
    if (arc_index == 1942) return "E"  ;
    if (arc_index == 1956) return "E"  ;
    if (arc_index == 2162) return "E"  ;
    if (arc_index == 2173) return "H"  ;
    if (arc_index == 2230) return "H"  ;
    if (arc_index == 2328) return "H"  ;
    if (arc_index == 2461) return "H"  ;
    if (arc_index == 2469) return "H"  ;
    if (arc_index == 2515) return "W"  ;
    if (arc_index == 2552) return "W"  ;
    if (arc_index == 2556) return "H"  ;
    if (arc_index == 2574) return "H"  ;
    if (arc_index == 2576) return "H"  ;
    if (arc_index == 2579) return "H"  ;
    if (arc_index == 2580) return "H"  ;
    if (arc_index == 2581) return "W"  ;
    if (arc_index == 2582) return "W"  ;
    if (arc_index == 2583) return "W"  ;
    if (arc_index == 2585) return "W"  ;
    if (arc_index == 2589) return "W"  ;
    if (arc_index == 2590) return "W"  ;
    if (arc_index == 2593) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2682) return "H"  ;
    if (arc_index == 2793) return "H"  ;
    if (arc_index == 2811) return "H"  ;
    if (arc_index == 2851) return "H"  ;
    if (arc_index == 2863) return "H"  ;
    if (arc_index == 2879) return "E"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 5)) begin 
    if (arc_index == 27) return "E"  ;
    if (arc_index == 134) return "H"  ;
    if (arc_index == 137) return "H"  ;
    if (arc_index == 139) return "E"  ;
    if (arc_index == 140) return "E"  ;
    if (arc_index == 143) return "E"  ;
    if (arc_index == 146) return "E"  ;
    if (arc_index == 147) return "E"  ;
    if (arc_index == 150) return "E"  ;
    if (arc_index == 223) return "W"  ;
    if (arc_index == 331) return "H"  ;
    if (arc_index == 374) return "H"  ;
    if (arc_index == 396) return "E"  ;
    if (arc_index == 397) return "E"  ;
    if (arc_index == 398) return "W"  ;
    if (arc_index == 399) return "W"  ;
    if (arc_index == 400) return "W"  ;
    if (arc_index == 401) return "W"  ;
    if (arc_index == 402) return "W"  ;
    if (arc_index == 403) return "W"  ;
    if (arc_index == 404) return "W"  ;
    if (arc_index == 405) return "W"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 407) return "W"  ;
    if (arc_index == 408) return "W"  ;
    if (arc_index == 409) return "W"  ;
    if (arc_index == 410) return "W"  ;
    if (arc_index == 411) return "W"  ;
    if (arc_index == 412) return "W"  ;
    if (arc_index == 413) return "W"  ;
    if (arc_index == 414) return "W"  ;
    if (arc_index == 415) return "W"  ;
    if (arc_index == 416) return "E"  ;
    if (arc_index == 417) return "W"  ;
    if (arc_index == 429) return "H"  ;
    if (arc_index == 474) return "H"  ;
    if (arc_index == 595) return "W"  ;
    if (arc_index == 660) return "W"  ;
    if (arc_index == 661) return "E"  ;
    if (arc_index == 671) return "E"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 673) return "H"  ;
    if (arc_index == 677) return "H"  ;
    if (arc_index == 680) return "E"  ;
    if (arc_index == 727) return "W"  ;
    if (arc_index == 728) return "W"  ;
    if (arc_index == 732) return "W"  ;
    if (arc_index == 738) return "W"  ;
    if (arc_index == 793) return "E"  ;
    if (arc_index == 804) return "E"  ;
    if (arc_index == 850) return "H"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 859) return "W"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 870) return "W"  ;
    if (arc_index == 875) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 878) return "W"  ;
    if (arc_index == 934) return "H"  ;
    if (arc_index == 936) return "E"  ;
    if (arc_index == 984) return "W"  ;
    if (arc_index == 1012) return "W"  ;
    if (arc_index == 1043) return "H"  ;
    if (arc_index == 1114) return "W"  ;
    if (arc_index == 1129) return "W"  ;
    if (arc_index == 1159) return "H"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1171) return "W"  ;
    if (arc_index == 1248) return "H"  ;
    if (arc_index == 1258) return "W"  ;
    if (arc_index == 1262) return "H"  ;
    if (arc_index == 1307) return "W"  ;
    if (arc_index == 1371) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1378) return "W"  ;
    if (arc_index == 1381) return "W"  ;
    if (arc_index == 1384) return "W"  ;
    if (arc_index == 1393) return "H"  ;
    if (arc_index == 1512) return "W"  ;
    if (arc_index == 1513) return "E"  ;
    if (arc_index == 1546) return "H"  ;
    if (arc_index == 1565) return "W"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1710) return "E"  ;
    if (arc_index == 1724) return "E"  ;
    if (arc_index == 1810) return "W"  ;
    if (arc_index == 1855) return "E"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2008) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2011) return "E"  ;
    if (arc_index == 2016) return "E"  ;
    if (arc_index == 2018) return "E"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2086) return "W"  ;
    if (arc_index == 2195) return "H"  ;
    if (arc_index == 2219) return "W"  ;
    if (arc_index == 2230) return "E"  ;
    if (arc_index == 2314) return "W"  ;
    if (arc_index == 2350) return "H"  ;
    if (arc_index == 2483) return "H"  ;
    if (arc_index == 2491) return "H"  ;
    if (arc_index == 2514) return "E"  ;
    if (arc_index == 2578) return "H"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2704) return "H"  ;
    if (arc_index == 2812) return "E"  ;
    if (arc_index == 2815) return "H"  ;
    if (arc_index == 2885) return "H"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 7)) begin 
    if (arc_index == 37) return "E"  ;
    if (arc_index == 90) return "W"  ;
    if (arc_index == 108) return "W"  ;
    if (arc_index == 126) return "E"  ;
    if (arc_index == 139) return "E"  ;
    if (arc_index == 140) return "E"  ;
    if (arc_index == 146) return "E"  ;
    if (arc_index == 147) return "E"  ;
    if (arc_index == 150) return "E"  ;
    if (arc_index == 156) return "H"  ;
    if (arc_index == 237) return "H"  ;
    if (arc_index == 287) return "W"  ;
    if (arc_index == 353) return "H"  ;
    if (arc_index == 354) return "H"  ;
    if (arc_index == 361) return "E"  ;
    if (arc_index == 364) return "E"  ;
    if (arc_index == 365) return "E"  ;
    if (arc_index == 370) return "E"  ;
    if (arc_index == 396) return "H"  ;
    if (arc_index == 416) return "E"  ;
    if (arc_index == 418) return "W"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 420) return "W"  ;
    if (arc_index == 421) return "W"  ;
    if (arc_index == 422) return "W"  ;
    if (arc_index == 423) return "E"  ;
    if (arc_index == 424) return "E"  ;
    if (arc_index == 425) return "E"  ;
    if (arc_index == 426) return "E"  ;
    if (arc_index == 427) return "E"  ;
    if (arc_index == 428) return "E"  ;
    if (arc_index == 429) return "W"  ;
    if (arc_index == 430) return "W"  ;
    if (arc_index == 431) return "W"  ;
    if (arc_index == 432) return "E"  ;
    if (arc_index == 433) return "E"  ;
    if (arc_index == 434) return "W"  ;
    if (arc_index == 435) return "E"  ;
    if (arc_index == 436) return "E"  ;
    if (arc_index == 437) return "E"  ;
    if (arc_index == 438) return "E"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 451) return "H"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 496) return "H"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 533) return "E"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 695) return "H"  ;
    if (arc_index == 735) return "H"  ;
    if (arc_index == 825) return "W"  ;
    if (arc_index == 857) return "W"  ;
    if (arc_index == 872) return "H"  ;
    if (arc_index == 944) return "H"  ;
    if (arc_index == 956) return "H"  ;
    if (arc_index == 1003) return "H"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1041) return "W"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1046) return "W"  ;
    if (arc_index == 1065) return "H"  ;
    if (arc_index == 1102) return "H"  ;
    if (arc_index == 1123) return "W"  ;
    if (arc_index == 1129) return "W"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1139) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1180) return "W"  ;
    if (arc_index == 1181) return "H"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1234) return "W"  ;
    if (arc_index == 1258) return "W"  ;
    if (arc_index == 1270) return "H"  ;
    if (arc_index == 1284) return "H"  ;
    if (arc_index == 1299) return "H"  ;
    if (arc_index == 1308) return "H"  ;
    if (arc_index == 1312) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1315) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1365) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1367) return "W"  ;
    if (arc_index == 1368) return "W"  ;
    if (arc_index == 1370) return "W"  ;
    if (arc_index == 1374) return "W"  ;
    if (arc_index == 1375) return "W"  ;
    if (arc_index == 1376) return "E"  ;
    if (arc_index == 1377) return "E"  ;
    if (arc_index == 1379) return "E"  ;
    if (arc_index == 1380) return "E"  ;
    if (arc_index == 1382) return "E"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1385) return "W"  ;
    if (arc_index == 1397) return "W"  ;
    if (arc_index == 1415) return "H"  ;
    if (arc_index == 1442) return "H"  ;
    if (arc_index == 1456) return "E"  ;
    if (arc_index == 1497) return "E"  ;
    if (arc_index == 1501) return "E"  ;
    if (arc_index == 1510) return "E"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1568) return "H"  ;
    if (arc_index == 1569) return "H"  ;
    if (arc_index == 1571) return "H"  ;
    if (arc_index == 1574) return "W"  ;
    if (arc_index == 1640) return "W"  ;
    if (arc_index == 1641) return "W"  ;
    if (arc_index == 1723) return "W"  ;
    if (arc_index == 1818) return "W"  ;
    if (arc_index == 1902) return "W"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1988) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2017) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2061) return "E"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2086) return "W"  ;
    if (arc_index == 2119) return "E"  ;
    if (arc_index == 2127) return "E"  ;
    if (arc_index == 2135) return "E"  ;
    if (arc_index == 2150) return "E"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2180) return "W"  ;
    if (arc_index == 2195) return "W"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2204) return "W"  ;
    if (arc_index == 2212) return "W"  ;
    if (arc_index == 2216) return "W"  ;
    if (arc_index == 2217) return "H"  ;
    if (arc_index == 2219) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2314) return "E"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2361) return "W"  ;
    if (arc_index == 2372) return "H"  ;
    if (arc_index == 2377) return "W"  ;
    if (arc_index == 2444) return "W"  ;
    if (arc_index == 2448) return "E"  ;
    if (arc_index == 2455) return "E"  ;
    if (arc_index == 2462) return "E"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2505) return "H"  ;
    if (arc_index == 2513) return "H"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2577) return "E"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2600) return "H"  ;
    if (arc_index == 2646) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2660) return "W"  ;
    if (arc_index == 2726) return "H"  ;
    if (arc_index == 2813) return "H"  ;
    if (arc_index == 2837) return "H"  ;
    if (arc_index == 2907) return "H"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 1)) begin 
    if (arc_index == 3) return "H"  ;
    if (arc_index == 47) return "W"  ;
    if (arc_index == 59) return "W"  ;
    if (arc_index == 69) return "W"  ;
    if (arc_index == 83) return "W"  ;
    if (arc_index == 145) return "W"  ;
    if (arc_index == 178) return "H"  ;
    if (arc_index == 222) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 375) return "H"  ;
    if (arc_index == 380) return "E"  ;
    if (arc_index == 384) return "E"  ;
    if (arc_index == 388) return "E"  ;
    if (arc_index == 389) return "E"  ;
    if (arc_index == 390) return "E"  ;
    if (arc_index == 395) return "E"  ;
    if (arc_index == 418) return "H"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 440) return "W"  ;
    if (arc_index == 441) return "W"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 443) return "E"  ;
    if (arc_index == 444) return "E"  ;
    if (arc_index == 445) return "E"  ;
    if (arc_index == 446) return "E"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 448) return "E"  ;
    if (arc_index == 449) return "E"  ;
    if (arc_index == 450) return "E"  ;
    if (arc_index == 451) return "E"  ;
    if (arc_index == 452) return "E"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 454) return "E"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 456) return "E"  ;
    if (arc_index == 457) return "W"  ;
    if (arc_index == 458) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 460) return "E"  ;
    if (arc_index == 461) return "E"  ;
    if (arc_index == 462) return "W"  ;
    if (arc_index == 473) return "H"  ;
    if (arc_index == 484) return "H"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 490) return "E"  ;
    if (arc_index == 495) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 497) return "E"  ;
    if (arc_index == 498) return "E"  ;
    if (arc_index == 501) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 513) return "E"  ;
    if (arc_index == 514) return "E"  ;
    if (arc_index == 517) return "W"  ;
    if (arc_index == 518) return "H"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 579) return "E"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 582) return "E"  ;
    if (arc_index == 592) return "E"  ;
    if (arc_index == 641) return "E"  ;
    if (arc_index == 717) return "H"  ;
    if (arc_index == 773) return "H"  ;
    if (arc_index == 800) return "H"  ;
    if (arc_index == 809) return "H"  ;
    if (arc_index == 894) return "H"  ;
    if (arc_index == 912) return "H"  ;
    if (arc_index == 924) return "H"  ;
    if (arc_index == 938) return "W"  ;
    if (arc_index == 948) return "W"  ;
    if (arc_index == 957) return "E"  ;
    if (arc_index == 978) return "H"  ;
    if (arc_index == 979) return "H"  ;
    if (arc_index == 1013) return "H"  ;
    if (arc_index == 1017) return "H"  ;
    if (arc_index == 1018) return "H"  ;
    if (arc_index == 1024) return "H"  ;
    if (arc_index == 1026) return "W"  ;
    if (arc_index == 1029) return "E"  ;
    if (arc_index == 1087) return "H"  ;
    if (arc_index == 1090) return "H"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1203) return "H"  ;
    if (arc_index == 1213) return "H"  ;
    if (arc_index == 1216) return "E"  ;
    if (arc_index == 1219) return "W"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1223) return "E"  ;
    if (arc_index == 1224) return "E"  ;
    if (arc_index == 1225) return "E"  ;
    if (arc_index == 1231) return "E"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1292) return "H"  ;
    if (arc_index == 1306) return "H"  ;
    if (arc_index == 1318) return "H"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1437) return "H"  ;
    if (arc_index == 1499) return "H"  ;
    if (arc_index == 1527) return "H"  ;
    if (arc_index == 1538) return "E"  ;
    if (arc_index == 1590) return "H"  ;
    if (arc_index == 1634) return "W"  ;
    if (arc_index == 1659) return "W"  ;
    if (arc_index == 1664) return "W"  ;
    if (arc_index == 1748) return "W"  ;
    if (arc_index == 1830) return "W"  ;
    if (arc_index == 1937) return "E"  ;
    if (arc_index == 1942) return "E"  ;
    if (arc_index == 1951) return "E"  ;
    if (arc_index == 1956) return "E"  ;
    if (arc_index == 2014) return "E"  ;
    if (arc_index == 2021) return "E"  ;
    if (arc_index == 2165) return "W"  ;
    if (arc_index == 2173) return "W"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2226) return "E"  ;
    if (arc_index == 2230) return "E"  ;
    if (arc_index == 2234) return "E"  ;
    if (arc_index == 2239) return "H"  ;
    if (arc_index == 2283) return "W"  ;
    if (arc_index == 2394) return "H"  ;
    if (arc_index == 2423) return "H"  ;
    if (arc_index == 2438) return "W"  ;
    if (arc_index == 2469) return "W"  ;
    if (arc_index == 2527) return "H"  ;
    if (arc_index == 2535) return "H"  ;
    if (arc_index == 2552) return "H"  ;
    if (arc_index == 2556) return "H"  ;
    if (arc_index == 2574) return "H"  ;
    if (arc_index == 2576) return "H"  ;
    if (arc_index == 2579) return "W"  ;
    if (arc_index == 2580) return "E"  ;
    if (arc_index == 2582) return "E"  ;
    if (arc_index == 2583) return "E"  ;
    if (arc_index == 2585) return "E"  ;
    if (arc_index == 2590) return "E"  ;
    if (arc_index == 2593) return "E"  ;
    if (arc_index == 2607) return "E"  ;
    if (arc_index == 2622) return "H"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2672) return "E"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2682) return "E"  ;
    if (arc_index == 2747) return "E"  ;
    if (arc_index == 2748) return "H"  ;
    if (arc_index == 2811) return "H"  ;
    if (arc_index == 2851) return "H"  ;
    if (arc_index == 2859) return "H"  ;
    if (arc_index == 2863) return "H"  ;
    if (arc_index == 2874) return "H"  ;
    if (arc_index == 2878) return "H"  ;
    if (arc_index == 2879) return "H"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 3)) begin 
    if (arc_index == 13) return "W"  ;
    if (arc_index == 18) return "W"  ;
    if (arc_index == 25) return "H"  ;
    if (arc_index == 35) return "H"  ;
    if (arc_index == 41) return "H"  ;
    if (arc_index == 49) return "H"  ;
    if (arc_index == 50) return "H"  ;
    if (arc_index == 63) return "W"  ;
    if (arc_index == 65) return "W"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 78) return "E"  ;
    if (arc_index == 81) return "E"  ;
    if (arc_index == 84) return "E"  ;
    if (arc_index == 86) return "E"  ;
    if (arc_index == 148) return "W"  ;
    if (arc_index == 152) return "W"  ;
    if (arc_index == 158) return "W"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 200) return "H"  ;
    if (arc_index == 216) return "H"  ;
    if (arc_index == 246) return "H"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 284) return "W"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 397) return "H"  ;
    if (arc_index == 404) return "H"  ;
    if (arc_index == 405) return "H"  ;
    if (arc_index == 406) return "H"  ;
    if (arc_index == 440) return "H"  ;
    if (arc_index == 454) return "H"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 456) return "E"  ;
    if (arc_index == 462) return "W"  ;
    if (arc_index == 463) return "E"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 465) return "W"  ;
    if (arc_index == 466) return "W"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 468) return "E"  ;
    if (arc_index == 469) return "E"  ;
    if (arc_index == 470) return "E"  ;
    if (arc_index == 471) return "E"  ;
    if (arc_index == 472) return "E"  ;
    if (arc_index == 473) return "W"  ;
    if (arc_index == 474) return "E"  ;
    if (arc_index == 475) return "E"  ;
    if (arc_index == 476) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 478) return "E"  ;
    if (arc_index == 479) return "E"  ;
    if (arc_index == 480) return "E"  ;
    if (arc_index == 481) return "E"  ;
    if (arc_index == 482) return "E"  ;
    if (arc_index == 483) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 495) return "H"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 540) return "H"  ;
    if (arc_index == 553) return "H"  ;
    if (arc_index == 562) return "H"  ;
    if (arc_index == 570) return "H"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 664) return "W"  ;
    if (arc_index == 668) return "W"  ;
    if (arc_index == 675) return "W"  ;
    if (arc_index == 676) return "W"  ;
    if (arc_index == 678) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 693) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 739) return "H"  ;
    if (arc_index == 750) return "H"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 811) return "E"  ;
    if (arc_index == 837) return "W"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 888) return "E"  ;
    if (arc_index == 895) return "E"  ;
    if (arc_index == 903) return "E"  ;
    if (arc_index == 904) return "E"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 910) return "E"  ;
    if (arc_index == 911) return "E"  ;
    if (arc_index == 914) return "E"  ;
    if (arc_index == 916) return "H"  ;
    if (arc_index == 917) return "E"  ;
    if (arc_index == 919) return "E"  ;
    if (arc_index == 920) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 923) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 980) return "W"  ;
    if (arc_index == 987) return "W"  ;
    if (arc_index == 994) return "W"  ;
    if (arc_index == 995) return "W"  ;
    if (arc_index == 1000) return "H"  ;
    if (arc_index == 1004) return "H"  ;
    if (arc_index == 1016) return "H"  ;
    if (arc_index == 1017) return "E"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1032) return "E"  ;
    if (arc_index == 1063) return "W"  ;
    if (arc_index == 1068) return "W"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1109) return "H"  ;
    if (arc_index == 1143) return "H"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1190) return "W"  ;
    if (arc_index == 1197) return "E"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1225) return "H"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1314) return "H"  ;
    if (arc_index == 1328) return "H"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1438) return "W"  ;
    if (arc_index == 1440) return "W"  ;
    if (arc_index == 1459) return "H"  ;
    if (arc_index == 1495) return "H"  ;
    if (arc_index == 1539) return "E"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1605) return "E"  ;
    if (arc_index == 1612) return "H"  ;
    if (arc_index == 1631) return "H"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1649) return "E"  ;
    if (arc_index == 1657) return "E"  ;
    if (arc_index == 1658) return "E"  ;
    if (arc_index == 1659) return "E"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1669) return "E"  ;
    if (arc_index == 1676) return "E"  ;
    if (arc_index == 1683) return "E"  ;
    if (arc_index == 1690) return "W"  ;
    if (arc_index == 1715) return "W"  ;
    if (arc_index == 1724) return "W"  ;
    if (arc_index == 1753) return "W"  ;
    if (arc_index == 1785) return "W"  ;
    if (arc_index == 1789) return "W"  ;
    if (arc_index == 1790) return "W"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1823) return "W"  ;
    if (arc_index == 1834) return "E"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1842) return "E"  ;
    if (arc_index == 1843) return "E"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1899) return "W"  ;
    if (arc_index == 1913) return "W"  ;
    if (arc_index == 1931) return "W"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1949) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 1960) return "W"  ;
    if (arc_index == 1987) return "W"  ;
    if (arc_index == 2001) return "W"  ;
    if (arc_index == 2013) return "W"  ;
    if (arc_index == 2023) return "W"  ;
    if (arc_index == 2024) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2035) return "W"  ;
    if (arc_index == 2040) return "W"  ;
    if (arc_index == 2052) return "W"  ;
    if (arc_index == 2066) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2116) return "W"  ;
    if (arc_index == 2155) return "W"  ;
    if (arc_index == 2157) return "W"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2166) return "W"  ;
    if (arc_index == 2170) return "W"  ;
    if (arc_index == 2171) return "W"  ;
    if (arc_index == 2172) return "E"  ;
    if (arc_index == 2176) return "W"  ;
    if (arc_index == 2177) return "W"  ;
    if (arc_index == 2222) return "E"  ;
    if (arc_index == 2227) return "E"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2235) return "E"  ;
    if (arc_index == 2236) return "E"  ;
    if (arc_index == 2237) return "E"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2243) return "E"  ;
    if (arc_index == 2248) return "W"  ;
    if (arc_index == 2255) return "W"  ;
    if (arc_index == 2261) return "H"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2416) return "H"  ;
    if (arc_index == 2421) return "H"  ;
    if (arc_index == 2422) return "H"  ;
    if (arc_index == 2429) return "E"  ;
    if (arc_index == 2432) return "E"  ;
    if (arc_index == 2434) return "E"  ;
    if (arc_index == 2442) return "E"  ;
    if (arc_index == 2450) return "W"  ;
    if (arc_index == 2460) return "W"  ;
    if (arc_index == 2475) return "E"  ;
    if (arc_index == 2483) return "E"  ;
    if (arc_index == 2485) return "W"  ;
    if (arc_index == 2486) return "W"  ;
    if (arc_index == 2508) return "W"  ;
    if (arc_index == 2516) return "W"  ;
    if (arc_index == 2535) return "W"  ;
    if (arc_index == 2540) return "W"  ;
    if (arc_index == 2549) return "H"  ;
    if (arc_index == 2557) return "H"  ;
    if (arc_index == 2566) return "E"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2589) return "E"  ;
    if (arc_index == 2644) return "H"  ;
    if (arc_index == 2662) return "H"  ;
    if (arc_index == 2664) return "E"  ;
    if (arc_index == 2669) return "E"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2694) return "E"  ;
    if (arc_index == 2697) return "E"  ;
    if (arc_index == 2704) return "E"  ;
    if (arc_index == 2713) return "E"  ;
    if (arc_index == 2755) return "E"  ;
    if (arc_index == 2770) return "H"  ;
    if (arc_index == 2793) return "H"  ;
    if (arc_index == 2796) return "H"  ;
    if (arc_index == 2803) return "H"  ;
    if (arc_index == 2842) return "H"  ;
    if (arc_index == 2854) return "H"  ;
    if (arc_index == 2856) return "W"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2881) return "H"  ;
    if (arc_index == 2887) return "H"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 0)) begin 
    if (arc_index == 47) return "H"  ;
    if (arc_index == 135) return "H"  ;
    if (arc_index == 222) return "H"  ;
    if (arc_index == 383) return "H"  ;
    if (arc_index == 419) return "H"  ;
    if (arc_index == 457) return "H"  ;
    if (arc_index == 462) return "H"  ;
    if (arc_index == 484) return "E"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 486) return "E"  ;
    if (arc_index == 487) return "E"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 490) return "E"  ;
    if (arc_index == 491) return "E"  ;
    if (arc_index == 492) return "E"  ;
    if (arc_index == 493) return "E"  ;
    if (arc_index == 494) return "E"  ;
    if (arc_index == 495) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 497) return "E"  ;
    if (arc_index == 498) return "E"  ;
    if (arc_index == 499) return "E"  ;
    if (arc_index == 500) return "E"  ;
    if (arc_index == 501) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 505) return "E"  ;
    if (arc_index == 517) return "H"  ;
    if (arc_index == 562) return "H"  ;
    if (arc_index == 575) return "H"  ;
    if (arc_index == 579) return "E"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 592) return "E"  ;
    if (arc_index == 761) return "H"  ;
    if (arc_index == 774) return "H"  ;
    if (arc_index == 938) return "H"  ;
    if (arc_index == 947) return "H"  ;
    if (arc_index == 1022) return "H"  ;
    if (arc_index == 1026) return "H"  ;
    if (arc_index == 1081) return "H"  ;
    if (arc_index == 1131) return "H"  ;
    if (arc_index == 1219) return "H"  ;
    if (arc_index == 1247) return "H"  ;
    if (arc_index == 1336) return "H"  ;
    if (arc_index == 1350) return "H"  ;
    if (arc_index == 1453) return "H"  ;
    if (arc_index == 1481) return "H"  ;
    if (arc_index == 1519) return "H"  ;
    if (arc_index == 1527) return "E"  ;
    if (arc_index == 1532) return "E"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1535) return "E"  ;
    if (arc_index == 1538) return "E"  ;
    if (arc_index == 1562) return "E"  ;
    if (arc_index == 1589) return "E"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1596) return "E"  ;
    if (arc_index == 1602) return "E"  ;
    if (arc_index == 1603) return "E"  ;
    if (arc_index == 1634) return "H"  ;
    if (arc_index == 2165) return "H"  ;
    if (arc_index == 2283) return "H"  ;
    if (arc_index == 2436) return "H"  ;
    if (arc_index == 2438) return "H"  ;
    if (arc_index == 2571) return "H"  ;
    if (arc_index == 2579) return "H"  ;
    if (arc_index == 2581) return "H"  ;
    if (arc_index == 2666) return "H"  ;
    if (arc_index == 2668) return "H"  ;
    if (arc_index == 2792) return "H"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2903) return "H"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 1)) begin 
    if (arc_index == 65) return "W"  ;
    if (arc_index == 69) return "H"  ;
    if (arc_index == 79) return "H"  ;
    if (arc_index == 106) return "H"  ;
    if (arc_index == 145) return "H"  ;
    if (arc_index == 244) return "H"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 389) return "W"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 441) return "H"  ;
    if (arc_index == 449) return "H"  ;
    if (arc_index == 450) return "H"  ;
    if (arc_index == 460) return "H"  ;
    if (arc_index == 478) return "H"  ;
    if (arc_index == 484) return "H"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 486) return "E"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 507) return "W"  ;
    if (arc_index == 508) return "W"  ;
    if (arc_index == 509) return "W"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 512) return "E"  ;
    if (arc_index == 513) return "E"  ;
    if (arc_index == 514) return "E"  ;
    if (arc_index == 515) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 517) return "E"  ;
    if (arc_index == 518) return "E"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 520) return "E"  ;
    if (arc_index == 521) return "E"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 523) return "E"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 539) return "H"  ;
    if (arc_index == 550) return "W"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 574) return "E"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 584) return "H"  ;
    if (arc_index == 589) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 591) return "E"  ;
    if (arc_index == 593) return "E"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 641) return "W"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 668) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 753) return "W"  ;
    if (arc_index == 773) return "W"  ;
    if (arc_index == 774) return "W"  ;
    if (arc_index == 783) return "H"  ;
    if (arc_index == 800) return "H"  ;
    if (arc_index == 840) return "W"  ;
    if (arc_index == 894) return "W"  ;
    if (arc_index == 924) return "W"  ;
    if (arc_index == 946) return "W"  ;
    if (arc_index == 948) return "W"  ;
    if (arc_index == 953) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 960) return "H"  ;
    if (arc_index == 962) return "H"  ;
    if (arc_index == 964) return "H"  ;
    if (arc_index == 965) return "E"  ;
    if (arc_index == 979) return "W"  ;
    if (arc_index == 1013) return "W"  ;
    if (arc_index == 1018) return "W"  ;
    if (arc_index == 1024) return "W"  ;
    if (arc_index == 1044) return "H"  ;
    if (arc_index == 1081) return "H"  ;
    if (arc_index == 1087) return "H"  ;
    if (arc_index == 1090) return "H"  ;
    if (arc_index == 1095) return "H"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1097) return "E"  ;
    if (arc_index == 1099) return "E"  ;
    if (arc_index == 1110) return "W"  ;
    if (arc_index == 1153) return "H"  ;
    if (arc_index == 1223) return "W"  ;
    if (arc_index == 1224) return "W"  ;
    if (arc_index == 1269) return "H"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1358) return "H"  ;
    if (arc_index == 1372) return "H"  ;
    if (arc_index == 1391) return "H"  ;
    if (arc_index == 1438) return "W"  ;
    if (arc_index == 1453) return "W"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1503) return "H"  ;
    if (arc_index == 1532) return "H"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1585) return "E"  ;
    if (arc_index == 1586) return "E"  ;
    if (arc_index == 1587) return "E"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1600) return "E"  ;
    if (arc_index == 1656) return "H"  ;
    if (arc_index == 1662) return "W"  ;
    if (arc_index == 1748) return "W"  ;
    if (arc_index == 1861) return "W"  ;
    if (arc_index == 1918) return "W"  ;
    if (arc_index == 1930) return "W"  ;
    if (arc_index == 1941) return "E"  ;
    if (arc_index == 1943) return "W"  ;
    if (arc_index == 1944) return "W"  ;
    if (arc_index == 1955) return "W"  ;
    if (arc_index == 1957) return "W"  ;
    if (arc_index == 2038) return "W"  ;
    if (arc_index == 2115) return "W"  ;
    if (arc_index == 2116) return "W"  ;
    if (arc_index == 2176) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2228) return "W"  ;
    if (arc_index == 2232) return "W"  ;
    if (arc_index == 2242) return "W"  ;
    if (arc_index == 2305) return "H"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2460) return "H"  ;
    if (arc_index == 2474) return "H"  ;
    if (arc_index == 2499) return "H"  ;
    if (arc_index == 2526) return "W"  ;
    if (arc_index == 2552) return "W"  ;
    if (arc_index == 2555) return "E"  ;
    if (arc_index == 2556) return "E"  ;
    if (arc_index == 2561) return "E"  ;
    if (arc_index == 2566) return "E"  ;
    if (arc_index == 2571) return "E"  ;
    if (arc_index == 2585) return "E"  ;
    if (arc_index == 2593) return "H"  ;
    if (arc_index == 2601) return "H"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2678) return "E"  ;
    if (arc_index == 2679) return "E"  ;
    if (arc_index == 2688) return "H"  ;
    if (arc_index == 2730) return "H"  ;
    if (arc_index == 2733) return "E"  ;
    if (arc_index == 2746) return "E"  ;
    if (arc_index == 2747) return "E"  ;
    if (arc_index == 2748) return "E"  ;
    if (arc_index == 2754) return "W"  ;
    if (arc_index == 2760) return "W"  ;
    if (arc_index == 2792) return "W"  ;
    if (arc_index == 2796) return "W"  ;
    if (arc_index == 2802) return "W"  ;
    if (arc_index == 2811) return "W"  ;
    if (arc_index == 2812) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2814) return "H"  ;
    if (arc_index == 2851) return "H"  ;
    if (arc_index == 2859) return "H"  ;
    if (arc_index == 2860) return "H"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2868) return "E"  ;
    if (arc_index == 2869) return "E"  ;
    if (arc_index == 2881) return "E"  ;
    if (arc_index == 2925) return "H"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 9)) begin 
    if (arc_index == 8) return "H"  ;
    if (arc_index == 21) return "H"  ;
    if (arc_index == 53) return "H"  ;
    if (arc_index == 56) return "H"  ;
    if (arc_index == 57) return "E"  ;
    if (arc_index == 91) return "H"  ;
    if (arc_index == 118) return "E"  ;
    if (arc_index == 119) return "E"  ;
    if (arc_index == 177) return "E"  ;
    if (arc_index == 183) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 192) return "W"  ;
    if (arc_index == 193) return "W"  ;
    if (arc_index == 209) return "E"  ;
    if (arc_index == 221) return "E"  ;
    if (arc_index == 234) return "E"  ;
    if (arc_index == 235) return "E"  ;
    if (arc_index == 236) return "E"  ;
    if (arc_index == 249) return "E"  ;
    if (arc_index == 250) return "E"  ;
    if (arc_index == 266) return "H"  ;
    if (arc_index == 283) return "H"  ;
    if (arc_index == 287) return "H"  ;
    if (arc_index == 295) return "H"  ;
    if (arc_index == 298) return "W"  ;
    if (arc_index == 303) return "W"  ;
    if (arc_index == 326) return "W"  ;
    if (arc_index == 348) return "W"  ;
    if (arc_index == 364) return "W"  ;
    if (arc_index == 402) return "E"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 425) return "E"  ;
    if (arc_index == 432) return "E"  ;
    if (arc_index == 463) return "H"  ;
    if (arc_index == 506) return "H"  ;
    if (arc_index == 528) return "H"  ;
    if (arc_index == 529) return "H"  ;
    if (arc_index == 530) return "W"  ;
    if (arc_index == 531) return "W"  ;
    if (arc_index == 532) return "W"  ;
    if (arc_index == 533) return "W"  ;
    if (arc_index == 534) return "W"  ;
    if (arc_index == 535) return "W"  ;
    if (arc_index == 536) return "W"  ;
    if (arc_index == 537) return "W"  ;
    if (arc_index == 538) return "W"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 540) return "W"  ;
    if (arc_index == 541) return "W"  ;
    if (arc_index == 542) return "W"  ;
    if (arc_index == 543) return "E"  ;
    if (arc_index == 544) return "E"  ;
    if (arc_index == 545) return "E"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 547) return "W"  ;
    if (arc_index == 548) return "W"  ;
    if (arc_index == 549) return "W"  ;
    if (arc_index == 561) return "H"  ;
    if (arc_index == 596) return "W"  ;
    if (arc_index == 606) return "H"  ;
    if (arc_index == 616) return "W"  ;
    if (arc_index == 620) return "W"  ;
    if (arc_index == 636) return "W"  ;
    if (arc_index == 639) return "W"  ;
    if (arc_index == 685) return "W"  ;
    if (arc_index == 725) return "W"  ;
    if (arc_index == 737) return "W"  ;
    if (arc_index == 741) return "W"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 805) return "H"  ;
    if (arc_index == 817) return "W"  ;
    if (arc_index == 818) return "E"  ;
    if (arc_index == 823) return "E"  ;
    if (arc_index == 825) return "E"  ;
    if (arc_index == 871) return "E"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 982) return "H"  ;
    if (arc_index == 1033) return "H"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1053) return "W"  ;
    if (arc_index == 1066) return "H"  ;
    if (arc_index == 1112) return "E"  ;
    if (arc_index == 1124) return "W"  ;
    if (arc_index == 1130) return "W"  ;
    if (arc_index == 1133) return "W"  ;
    if (arc_index == 1134) return "W"  ;
    if (arc_index == 1136) return "W"  ;
    if (arc_index == 1142) return "W"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1175) return "H"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1235) return "W"  ;
    if (arc_index == 1239) return "W"  ;
    if (arc_index == 1242) return "W"  ;
    if (arc_index == 1251) return "W"  ;
    if (arc_index == 1253) return "W"  ;
    if (arc_index == 1268) return "W"  ;
    if (arc_index == 1271) return "W"  ;
    if (arc_index == 1278) return "W"  ;
    if (arc_index == 1283) return "W"  ;
    if (arc_index == 1291) return "H"  ;
    if (arc_index == 1298) return "H"  ;
    if (arc_index == 1304) return "H"  ;
    if (arc_index == 1305) return "H"  ;
    if (arc_index == 1313) return "H"  ;
    if (arc_index == 1316) return "H"  ;
    if (arc_index == 1324) return "E"  ;
    if (arc_index == 1331) return "E"  ;
    if (arc_index == 1338) return "E"  ;
    if (arc_index == 1342) return "E"  ;
    if (arc_index == 1361) return "W"  ;
    if (arc_index == 1380) return "H"  ;
    if (arc_index == 1382) return "H"  ;
    if (arc_index == 1394) return "H"  ;
    if (arc_index == 1399) return "E"  ;
    if (arc_index == 1434) return "E"  ;
    if (arc_index == 1446) return "E"  ;
    if (arc_index == 1450) return "E"  ;
    if (arc_index == 1479) return "E"  ;
    if (arc_index == 1488) return "E"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1525) return "H"  ;
    if (arc_index == 1567) return "H"  ;
    if (arc_index == 1580) return "H"  ;
    if (arc_index == 1583) return "H"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1678) return "H"  ;
    if (arc_index == 1686) return "H"  ;
    if (arc_index == 1692) return "H"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1770) return "E"  ;
    if (arc_index == 1797) return "E"  ;
    if (arc_index == 1809) return "E"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1867) return "E"  ;
    if (arc_index == 1875) return "E"  ;
    if (arc_index == 1880) return "E"  ;
    if (arc_index == 1891) return "E"  ;
    if (arc_index == 1916) return "E"  ;
    if (arc_index == 1962) return "E"  ;
    if (arc_index == 1974) return "E"  ;
    if (arc_index == 1975) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2046) return "E"  ;
    if (arc_index == 2048) return "E"  ;
    if (arc_index == 2068) return "E"  ;
    if (arc_index == 2070) return "E"  ;
    if (arc_index == 2072) return "E"  ;
    if (arc_index == 2079) return "W"  ;
    if (arc_index == 2098) return "W"  ;
    if (arc_index == 2100) return "E"  ;
    if (arc_index == 2113) return "E"  ;
    if (arc_index == 2136) return "E"  ;
    if (arc_index == 2141) return "E"  ;
    if (arc_index == 2156) return "E"  ;
    if (arc_index == 2179) return "W"  ;
    if (arc_index == 2183) return "W"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2186) return "W"  ;
    if (arc_index == 2188) return "W"  ;
    if (arc_index == 2189) return "W"  ;
    if (arc_index == 2190) return "W"  ;
    if (arc_index == 2193) return "W"  ;
    if (arc_index == 2245) return "W"  ;
    if (arc_index == 2256) return "E"  ;
    if (arc_index == 2269) return "E"  ;
    if (arc_index == 2271) return "E"  ;
    if (arc_index == 2288) return "E"  ;
    if (arc_index == 2295) return "E"  ;
    if (arc_index == 2310) return "E"  ;
    if (arc_index == 2313) return "E"  ;
    if (arc_index == 2315) return "W"  ;
    if (arc_index == 2317) return "W"  ;
    if (arc_index == 2320) return "W"  ;
    if (arc_index == 2322) return "W"  ;
    if (arc_index == 2326) return "W"  ;
    if (arc_index == 2327) return "H"  ;
    if (arc_index == 2329) return "H"  ;
    if (arc_index == 2331) return "H"  ;
    if (arc_index == 2343) return "H"  ;
    if (arc_index == 2377) return "H"  ;
    if (arc_index == 2404) return "W"  ;
    if (arc_index == 2408) return "W"  ;
    if (arc_index == 2411) return "W"  ;
    if (arc_index == 2414) return "W"  ;
    if (arc_index == 2417) return "W"  ;
    if (arc_index == 2418) return "W"  ;
    if (arc_index == 2431) return "W"  ;
    if (arc_index == 2482) return "H"  ;
    if (arc_index == 2594) return "H"  ;
    if (arc_index == 2615) return "H"  ;
    if (arc_index == 2623) return "H"  ;
    if (arc_index == 2633) return "W"  ;
    if (arc_index == 2638) return "W"  ;
    if (arc_index == 2639) return "W"  ;
    if (arc_index == 2643) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2706) return "E"  ;
    if (arc_index == 2707) return "E"  ;
    if (arc_index == 2708) return "W"  ;
    if (arc_index == 2709) return "W"  ;
    if (arc_index == 2710) return "H"  ;
    if (arc_index == 2713) return "H"  ;
    if (arc_index == 2714) return "H"  ;
    if (arc_index == 2717) return "H"  ;
    if (arc_index == 2720) return "W"  ;
    if (arc_index == 2721) return "W"  ;
    if (arc_index == 2722) return "W"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2831) return "E"  ;
    if (arc_index == 2836) return "H"  ;
    if (arc_index == 2848) return "H"  ;
    if (arc_index == 2905) return "W"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 7)) begin 
    if (arc_index == 43) return "H"  ;
    if (arc_index == 113) return "H"  ;
    if (arc_index == 281) return "W"  ;
    if (arc_index == 288) return "H"  ;
    if (arc_index == 485) return "H"  ;
    if (arc_index == 528) return "H"  ;
    if (arc_index == 550) return "W"  ;
    if (arc_index == 551) return "E"  ;
    if (arc_index == 552) return "E"  ;
    if (arc_index == 553) return "W"  ;
    if (arc_index == 554) return "W"  ;
    if (arc_index == 555) return "W"  ;
    if (arc_index == 556) return "E"  ;
    if (arc_index == 557) return "E"  ;
    if (arc_index == 558) return "E"  ;
    if (arc_index == 559) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 561) return "W"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 563) return "E"  ;
    if (arc_index == 564) return "E"  ;
    if (arc_index == 565) return "W"  ;
    if (arc_index == 566) return "E"  ;
    if (arc_index == 567) return "W"  ;
    if (arc_index == 568) return "E"  ;
    if (arc_index == 569) return "W"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 571) return "W"  ;
    if (arc_index == 583) return "H"  ;
    if (arc_index == 628) return "H"  ;
    if (arc_index == 712) return "W"  ;
    if (arc_index == 788) return "E"  ;
    if (arc_index == 827) return "H"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 1004) return "H"  ;
    if (arc_index == 1088) return "H"  ;
    if (arc_index == 1197) return "H"  ;
    if (arc_index == 1313) return "H"  ;
    if (arc_index == 1343) return "W"  ;
    if (arc_index == 1402) return "H"  ;
    if (arc_index == 1409) return "H"  ;
    if (arc_index == 1416) return "H"  ;
    if (arc_index == 1420) return "H"  ;
    if (arc_index == 1426) return "E"  ;
    if (arc_index == 1472) return "E"  ;
    if (arc_index == 1498) return "E"  ;
    if (arc_index == 1547) return "H"  ;
    if (arc_index == 1695) return "E"  ;
    if (arc_index == 1700) return "H"  ;
    if (arc_index == 1701) return "E"  ;
    if (arc_index == 1708) return "E"  ;
    if (arc_index == 1714) return "E"  ;
    if (arc_index == 1761) return "W"  ;
    if (arc_index == 1762) return "W"  ;
    if (arc_index == 1767) return "W"  ;
    if (arc_index == 1771) return "W"  ;
    if (arc_index == 1772) return "W"  ;
    if (arc_index == 1838) return "E"  ;
    if (arc_index == 2025) return "E"  ;
    if (arc_index == 2037) return "E"  ;
    if (arc_index == 2094) return "W"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2099) return "W"  ;
    if (arc_index == 2102) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2110) return "W"  ;
    if (arc_index == 2298) return "E"  ;
    if (arc_index == 2335) return "W"  ;
    if (arc_index == 2341) return "W"  ;
    if (arc_index == 2349) return "H"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2504) return "H"  ;
    if (arc_index == 2544) return "E"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2637) return "H"  ;
    if (arc_index == 2645) return "H"  ;
    if (arc_index == 2732) return "H"  ;
    if (arc_index == 2737) return "E"  ;
    if (arc_index == 2777) return "E"  ;
    if (arc_index == 2853) return "E"  ;
    if (arc_index == 2858) return "H"  ;
    if (arc_index == 2916) return "W"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 0)) begin 
    if (arc_index == 65) return "H"  ;
    if (arc_index == 135) return "H"  ;
    if (arc_index == 310) return "H"  ;
    if (arc_index == 388) return "H"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 492) return "E"  ;
    if (arc_index == 493) return "E"  ;
    if (arc_index == 507) return "H"  ;
    if (arc_index == 509) return "H"  ;
    if (arc_index == 550) return "H"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 574) return "E"  ;
    if (arc_index == 575) return "E"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 577) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 579) return "E"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 581) return "E"  ;
    if (arc_index == 582) return "E"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 584) return "E"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 587) return "E"  ;
    if (arc_index == 588) return "E"  ;
    if (arc_index == 589) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 591) return "E"  ;
    if (arc_index == 592) return "E"  ;
    if (arc_index == 593) return "E"  ;
    if (arc_index == 605) return "H"  ;
    if (arc_index == 650) return "H"  ;
    if (arc_index == 753) return "H"  ;
    if (arc_index == 761) return "H"  ;
    if (arc_index == 840) return "H"  ;
    if (arc_index == 849) return "H"  ;
    if (arc_index == 924) return "H"  ;
    if (arc_index == 947) return "H"  ;
    if (arc_index == 957) return "H"  ;
    if (arc_index == 960) return "E"  ;
    if (arc_index == 964) return "E"  ;
    if (arc_index == 966) return "E"  ;
    if (arc_index == 979) return "E"  ;
    if (arc_index == 1024) return "E"  ;
    if (arc_index == 1026) return "H"  ;
    if (arc_index == 1110) return "H"  ;
    if (arc_index == 1219) return "H"  ;
    if (arc_index == 1223) return "H"  ;
    if (arc_index == 1335) return "H"  ;
    if (arc_index == 1424) return "H"  ;
    if (arc_index == 1438) return "H"  ;
    if (arc_index == 1481) return "H"  ;
    if (arc_index == 1569) return "H"  ;
    if (arc_index == 1585) return "E"  ;
    if (arc_index == 1586) return "E"  ;
    if (arc_index == 1587) return "E"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1593) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1600) return "E"  ;
    if (arc_index == 1601) return "E"  ;
    if (arc_index == 1662) return "E"  ;
    if (arc_index == 1722) return "H"  ;
    if (arc_index == 1861) return "H"  ;
    if (arc_index == 1943) return "H"  ;
    if (arc_index == 2021) return "H"  ;
    if (arc_index == 2038) return "H"  ;
    if (arc_index == 2044) return "H"  ;
    if (arc_index == 2116) return "H"  ;
    if (arc_index == 2242) return "H"  ;
    if (arc_index == 2371) return "H"  ;
    if (arc_index == 2423) return "H"  ;
    if (arc_index == 2526) return "H"  ;
    if (arc_index == 2659) return "H"  ;
    if (arc_index == 2663) return "H"  ;
    if (arc_index == 2667) return "H"  ;
    if (arc_index == 2671) return "H"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2678) return "E"  ;
    if (arc_index == 2679) return "E"  ;
    if (arc_index == 2734) return "E"  ;
    if (arc_index == 2740) return "E"  ;
    if (arc_index == 2754) return "H"  ;
    if (arc_index == 2792) return "H"  ;
    if (arc_index == 2860) return "E"  ;
    if (arc_index == 2863) return "E"  ;
    if (arc_index == 2868) return "E"  ;
    if (arc_index == 2869) return "E"  ;
    if (arc_index == 2874) return "E"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2879) return "E"  ;
    if (arc_index == 2880) return "H"  ;
    if (arc_index == 2881) return "E"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 10)) begin 
    if (arc_index == 87) return "H"  ;
    if (arc_index == 97) return "E"  ;
    if (arc_index == 157) return "H"  ;
    if (arc_index == 179) return "H"  ;
    if (arc_index == 191) return "H"  ;
    if (arc_index == 197) return "H"  ;
    if (arc_index == 203) return "H"  ;
    if (arc_index == 213) return "E"  ;
    if (arc_index == 254) return "E"  ;
    if (arc_index == 286) return "E"  ;
    if (arc_index == 288) return "E"  ;
    if (arc_index == 294) return "E"  ;
    if (arc_index == 300) return "E"  ;
    if (arc_index == 301) return "W"  ;
    if (arc_index == 302) return "E"  ;
    if (arc_index == 305) return "E"  ;
    if (arc_index == 307) return "E"  ;
    if (arc_index == 316) return "E"  ;
    if (arc_index == 319) return "E"  ;
    if (arc_index == 324) return "W"  ;
    if (arc_index == 332) return "H"  ;
    if (arc_index == 339) return "H"  ;
    if (arc_index == 341) return "H"  ;
    if (arc_index == 370) return "H"  ;
    if (arc_index == 455) return "H"  ;
    if (arc_index == 529) return "H"  ;
    if (arc_index == 563) return "H"  ;
    if (arc_index == 566) return "H"  ;
    if (arc_index == 572) return "H"  ;
    if (arc_index == 594) return "H"  ;
    if (arc_index == 595) return "W"  ;
    if (arc_index == 596) return "W"  ;
    if (arc_index == 597) return "W"  ;
    if (arc_index == 598) return "W"  ;
    if (arc_index == 599) return "W"  ;
    if (arc_index == 600) return "E"  ;
    if (arc_index == 601) return "E"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 603) return "W"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 606) return "W"  ;
    if (arc_index == 607) return "W"  ;
    if (arc_index == 608) return "W"  ;
    if (arc_index == 609) return "W"  ;
    if (arc_index == 610) return "W"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 613) return "W"  ;
    if (arc_index == 614) return "W"  ;
    if (arc_index == 615) return "W"  ;
    if (arc_index == 616) return "W"  ;
    if (arc_index == 620) return "W"  ;
    if (arc_index == 622) return "W"  ;
    if (arc_index == 627) return "H"  ;
    if (arc_index == 636) return "H"  ;
    if (arc_index == 639) return "H"  ;
    if (arc_index == 672) return "H"  ;
    if (arc_index == 701) return "H"  ;
    if (arc_index == 704) return "W"  ;
    if (arc_index == 714) return "W"  ;
    if (arc_index == 723) return "W"  ;
    if (arc_index == 725) return "W"  ;
    if (arc_index == 737) return "W"  ;
    if (arc_index == 741) return "W"  ;
    if (arc_index == 824) return "W"  ;
    if (arc_index == 871) return "H"  ;
    if (arc_index == 1034) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1048) return "H"  ;
    if (arc_index == 1050) return "H"  ;
    if (arc_index == 1067) return "H"  ;
    if (arc_index == 1071) return "H"  ;
    if (arc_index == 1122) return "H"  ;
    if (arc_index == 1132) return "H"  ;
    if (arc_index == 1141) return "H"  ;
    if (arc_index == 1152) return "H"  ;
    if (arc_index == 1155) return "H"  ;
    if (arc_index == 1163) return "H"  ;
    if (arc_index == 1241) return "H"  ;
    if (arc_index == 1242) return "H"  ;
    if (arc_index == 1277) return "H"  ;
    if (arc_index == 1305) return "H"  ;
    if (arc_index == 1320) return "H"  ;
    if (arc_index == 1326) return "H"  ;
    if (arc_index == 1339) return "H"  ;
    if (arc_index == 1342) return "H"  ;
    if (arc_index == 1347) return "H"  ;
    if (arc_index == 1354) return "W"  ;
    if (arc_index == 1357) return "H"  ;
    if (arc_index == 1361) return "H"  ;
    if (arc_index == 1446) return "H"  ;
    if (arc_index == 1460) return "H"  ;
    if (arc_index == 1475) return "H"  ;
    if (arc_index == 1544) return "W"  ;
    if (arc_index == 1554) return "W"  ;
    if (arc_index == 1570) return "W"  ;
    if (arc_index == 1577) return "W"  ;
    if (arc_index == 1591) return "H"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1744) return "H"  ;
    if (arc_index == 1769) return "H"  ;
    if (arc_index == 1806) return "H"  ;
    if (arc_index == 1869) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2081) return "W"  ;
    if (arc_index == 2089) return "W"  ;
    if (arc_index == 2101) return "W"  ;
    if (arc_index == 2181) return "W"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2194) return "W"  ;
    if (arc_index == 2196) return "W"  ;
    if (arc_index == 2198) return "W"  ;
    if (arc_index == 2208) return "W"  ;
    if (arc_index == 2303) return "W"  ;
    if (arc_index == 2345) return "W"  ;
    if (arc_index == 2354) return "E"  ;
    if (arc_index == 2373) return "E"  ;
    if (arc_index == 2376) return "E"  ;
    if (arc_index == 2377) return "E"  ;
    if (arc_index == 2381) return "E"  ;
    if (arc_index == 2382) return "E"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2386) return "W"  ;
    if (arc_index == 2387) return "W"  ;
    if (arc_index == 2389) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2393) return "H"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2395) return "W"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2537) return "E"  ;
    if (arc_index == 2548) return "H"  ;
    if (arc_index == 2623) return "H"  ;
    if (arc_index == 2632) return "H"  ;
    if (arc_index == 2633) return "H"  ;
    if (arc_index == 2638) return "H"  ;
    if (arc_index == 2639) return "H"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2681) return "H"  ;
    if (arc_index == 2689) return "H"  ;
    if (arc_index == 2690) return "H"  ;
    if (arc_index == 2696) return "H"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2727) return "W"  ;
    if (arc_index == 2776) return "H"  ;
    if (arc_index == 2825) return "H"  ;
    if (arc_index == 2830) return "E"  ;
    if (arc_index == 2833) return "E"  ;
    if (arc_index == 2895) return "E"  ;
    if (arc_index == 2902) return "H"  ;
    if (arc_index == 2905) return "H"  ;
    if (arc_index == 2907) return "W"  ;
    if (arc_index == 2913) return "W"  ;
    if (arc_index == 2920) return "W"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 11)) begin 
    if (arc_index == 109) return "H"  ;
    if (arc_index == 179) return "H"  ;
    if (arc_index == 354) return "H"  ;
    if (arc_index == 551) return "H"  ;
    if (arc_index == 558) return "H"  ;
    if (arc_index == 594) return "H"  ;
    if (arc_index == 616) return "H"  ;
    if (arc_index == 617) return "W"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 619) return "W"  ;
    if (arc_index == 620) return "W"  ;
    if (arc_index == 621) return "W"  ;
    if (arc_index == 622) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 625) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 627) return "W"  ;
    if (arc_index == 628) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 630) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 632) return "W"  ;
    if (arc_index == 633) return "W"  ;
    if (arc_index == 634) return "W"  ;
    if (arc_index == 635) return "W"  ;
    if (arc_index == 636) return "W"  ;
    if (arc_index == 637) return "W"  ;
    if (arc_index == 649) return "H"  ;
    if (arc_index == 694) return "H"  ;
    if (arc_index == 711) return "H"  ;
    if (arc_index == 893) return "H"  ;
    if (arc_index == 1070) return "H"  ;
    if (arc_index == 1154) return "H"  ;
    if (arc_index == 1263) return "H"  ;
    if (arc_index == 1379) return "H"  ;
    if (arc_index == 1468) return "H"  ;
    if (arc_index == 1482) return "H"  ;
    if (arc_index == 1556) return "W"  ;
    if (arc_index == 1613) return "H"  ;
    if (arc_index == 1766) return "H"  ;
    if (arc_index == 1777) return "H"  ;
    if (arc_index == 1779) return "H"  ;
    if (arc_index == 2111) return "H"  ;
    if (arc_index == 2415) return "H"  ;
    if (arc_index == 2570) return "H"  ;
    if (arc_index == 2626) return "W"  ;
    if (arc_index == 2628) return "W"  ;
    if (arc_index == 2629) return "W"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2635) return "W"  ;
    if (arc_index == 2636) return "W"  ;
    if (arc_index == 2637) return "W"  ;
    if (arc_index == 2658) return "W"  ;
    if (arc_index == 2703) return "H"  ;
    if (arc_index == 2711) return "H"  ;
    if (arc_index == 2798) return "H"  ;
    if (arc_index == 2906) return "W"  ;
    if (arc_index == 2910) return "W"  ;
    if (arc_index == 2916) return "W"  ;
    if (arc_index == 2923) return "W"  ;
    if (arc_index == 2924) return "H"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 6)) begin 
    if (arc_index == 19) return "H"  ;
    if (arc_index == 20) return "H"  ;
    if (arc_index == 23) return "E"  ;
    if (arc_index == 37) return "E"  ;
    if (arc_index == 66) return "E"  ;
    if (arc_index == 88) return "W"  ;
    if (arc_index == 93) return "W"  ;
    if (arc_index == 96) return "W"  ;
    if (arc_index == 98) return "W"  ;
    if (arc_index == 99) return "W"  ;
    if (arc_index == 100) return "W"  ;
    if (arc_index == 102) return "W"  ;
    if (arc_index == 106) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 111) return "E"  ;
    if (arc_index == 121) return "E"  ;
    if (arc_index == 126) return "E"  ;
    if (arc_index == 127) return "E"  ;
    if (arc_index == 131) return "H"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 188) return "W"  ;
    if (arc_index == 201) return "H"  ;
    if (arc_index == 223) return "H"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 330) return "W"  ;
    if (arc_index == 331) return "W"  ;
    if (arc_index == 351) return "W"  ;
    if (arc_index == 356) return "W"  ;
    if (arc_index == 358) return "W"  ;
    if (arc_index == 359) return "W"  ;
    if (arc_index == 362) return "W"  ;
    if (arc_index == 363) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 367) return "W"  ;
    if (arc_index == 371) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 376) return "H"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 385) return "E"  ;
    if (arc_index == 393) return "E"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 401) return "E"  ;
    if (arc_index == 402) return "E"  ;
    if (arc_index == 408) return "E"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 415) return "E"  ;
    if (arc_index == 426) return "E"  ;
    if (arc_index == 436) return "E"  ;
    if (arc_index == 451) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 564) return "W"  ;
    if (arc_index == 573) return "H"  ;
    if (arc_index == 595) return "H"  ;
    if (arc_index == 596) return "H"  ;
    if (arc_index == 616) return "H"  ;
    if (arc_index == 629) return "H"  ;
    if (arc_index == 638) return "H"  ;
    if (arc_index == 639) return "H"  ;
    if (arc_index == 640) return "W"  ;
    if (arc_index == 641) return "W"  ;
    if (arc_index == 642) return "W"  ;
    if (arc_index == 643) return "E"  ;
    if (arc_index == 644) return "W"  ;
    if (arc_index == 645) return "W"  ;
    if (arc_index == 646) return "E"  ;
    if (arc_index == 647) return "E"  ;
    if (arc_index == 648) return "W"  ;
    if (arc_index == 649) return "W"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 651) return "W"  ;
    if (arc_index == 652) return "E"  ;
    if (arc_index == 653) return "E"  ;
    if (arc_index == 654) return "E"  ;
    if (arc_index == 655) return "E"  ;
    if (arc_index == 656) return "E"  ;
    if (arc_index == 657) return "E"  ;
    if (arc_index == 658) return "E"  ;
    if (arc_index == 659) return "E"  ;
    if (arc_index == 660) return "E"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 671) return "H"  ;
    if (arc_index == 677) return "H"  ;
    if (arc_index == 716) return "H"  ;
    if (arc_index == 726) return "H"  ;
    if (arc_index == 744) return "H"  ;
    if (arc_index == 795) return "E"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 836) return "E"  ;
    if (arc_index == 863) return "E"  ;
    if (arc_index == 866) return "E"  ;
    if (arc_index == 868) return "E"  ;
    if (arc_index == 869) return "E"  ;
    if (arc_index == 876) return "E"  ;
    if (arc_index == 890) return "E"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 915) return "H"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 940) return "E"  ;
    if (arc_index == 941) return "E"  ;
    if (arc_index == 970) return "E"  ;
    if (arc_index == 992) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1069) return "E"  ;
    if (arc_index == 1085) return "E"  ;
    if (arc_index == 1092) return "H"  ;
    if (arc_index == 1102) return "E"  ;
    if (arc_index == 1107) return "W"  ;
    if (arc_index == 1114) return "W"  ;
    if (arc_index == 1115) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1171) return "W"  ;
    if (arc_index == 1176) return "H"  ;
    if (arc_index == 1180) return "H"  ;
    if (arc_index == 1181) return "H"  ;
    if (arc_index == 1189) return "E"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1218) return "E"  ;
    if (arc_index == 1240) return "W"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1245) return "W"  ;
    if (arc_index == 1246) return "W"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1260) return "W"  ;
    if (arc_index == 1262) return "W"  ;
    if (arc_index == 1267) return "W"  ;
    if (arc_index == 1272) return "W"  ;
    if (arc_index == 1282) return "W"  ;
    if (arc_index == 1285) return "H"  ;
    if (arc_index == 1303) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1365) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1368) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1396) return "W"  ;
    if (arc_index == 1401) return "H"  ;
    if (arc_index == 1442) return "E"  ;
    if (arc_index == 1456) return "E"  ;
    if (arc_index == 1474) return "W"  ;
    if (arc_index == 1490) return "H"  ;
    if (arc_index == 1504) return "H"  ;
    if (arc_index == 1509) return "E"  ;
    if (arc_index == 1555) return "E"  ;
    if (arc_index == 1563) return "E"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1621) return "W"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1635) return "H"  ;
    if (arc_index == 1640) return "H"  ;
    if (arc_index == 1677) return "W"  ;
    if (arc_index == 1687) return "W"  ;
    if (arc_index == 1764) return "W"  ;
    if (arc_index == 1788) return "H"  ;
    if (arc_index == 1810) return "H"  ;
    if (arc_index == 1878) return "W"  ;
    if (arc_index == 1890) return "W"  ;
    if (arc_index == 1902) return "E"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 2018) return "E"  ;
    if (arc_index == 2019) return "E"  ;
    if (arc_index == 2061) return "E"  ;
    if (arc_index == 2069) return "W"  ;
    if (arc_index == 2071) return "W"  ;
    if (arc_index == 2074) return "W"  ;
    if (arc_index == 2120) return "E"  ;
    if (arc_index == 2127) return "E"  ;
    if (arc_index == 2135) return "E"  ;
    if (arc_index == 2136) return "E"  ;
    if (arc_index == 2142) return "E"  ;
    if (arc_index == 2146) return "E"  ;
    if (arc_index == 2147) return "E"  ;
    if (arc_index == 2175) return "E"  ;
    if (arc_index == 2197) return "W"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2202) return "W"  ;
    if (arc_index == 2204) return "W"  ;
    if (arc_index == 2205) return "W"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2246) return "W"  ;
    if (arc_index == 2306) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2411) return "W"  ;
    if (arc_index == 2418) return "W"  ;
    if (arc_index == 2437) return "H"  ;
    if (arc_index == 2439) return "H"  ;
    if (arc_index == 2446) return "E"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2505) return "E"  ;
    if (arc_index == 2512) return "E"  ;
    if (arc_index == 2517) return "E"  ;
    if (arc_index == 2522) return "E"  ;
    if (arc_index == 2525) return "E"  ;
    if (arc_index == 2528) return "E"  ;
    if (arc_index == 2534) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2592) return "H"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2599) return "W"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2673) return "W"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2719) return "W"  ;
    if (arc_index == 2725) return "H"  ;
    if (arc_index == 2733) return "H"  ;
    if (arc_index == 2752) return "E"  ;
    if (arc_index == 2771) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2820) return "H"  ;
    if (arc_index == 2841) return "H"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 3)) begin 
    if (arc_index == 40) return "W"  ;
    if (arc_index == 42) return "H"  ;
    if (arc_index == 141) return "H"  ;
    if (arc_index == 144) return "H"  ;
    if (arc_index == 151) return "H"  ;
    if (arc_index == 153) return "H"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 223) return "H"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 398) return "H"  ;
    if (arc_index == 407) return "W"  ;
    if (arc_index == 411) return "W"  ;
    if (arc_index == 417) return "W"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 595) return "H"  ;
    if (arc_index == 638) return "H"  ;
    if (arc_index == 660) return "E"  ;
    if (arc_index == 661) return "E"  ;
    if (arc_index == 662) return "W"  ;
    if (arc_index == 663) return "W"  ;
    if (arc_index == 664) return "W"  ;
    if (arc_index == 665) return "E"  ;
    if (arc_index == 666) return "E"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 668) return "E"  ;
    if (arc_index == 669) return "E"  ;
    if (arc_index == 670) return "E"  ;
    if (arc_index == 671) return "E"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 673) return "E"  ;
    if (arc_index == 674) return "E"  ;
    if (arc_index == 675) return "E"  ;
    if (arc_index == 676) return "E"  ;
    if (arc_index == 677) return "E"  ;
    if (arc_index == 678) return "E"  ;
    if (arc_index == 679) return "E"  ;
    if (arc_index == 680) return "E"  ;
    if (arc_index == 681) return "W"  ;
    if (arc_index == 693) return "H"  ;
    if (arc_index == 738) return "H"  ;
    if (arc_index == 804) return "E"  ;
    if (arc_index == 859) return "W"  ;
    if (arc_index == 875) return "W"  ;
    if (arc_index == 934) return "E"  ;
    if (arc_index == 936) return "E"  ;
    if (arc_index == 937) return "H"  ;
    if (arc_index == 990) return "W"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1014) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1019) return "E"  ;
    if (arc_index == 1023) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1114) return "H"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1171) return "W"  ;
    if (arc_index == 1198) return "H"  ;
    if (arc_index == 1258) return "W"  ;
    if (arc_index == 1289) return "W"  ;
    if (arc_index == 1307) return "H"  ;
    if (arc_index == 1384) return "W"  ;
    if (arc_index == 1423) return "H"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1512) return "H"  ;
    if (arc_index == 1526) return "H"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1565) return "W"  ;
    if (arc_index == 1657) return "H"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1810) return "H"  ;
    if (arc_index == 1980) return "W"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2005) return "E"  ;
    if (arc_index == 2008) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2011) return "E"  ;
    if (arc_index == 2016) return "E"  ;
    if (arc_index == 2017) return "E"  ;
    if (arc_index == 2018) return "E"  ;
    if (arc_index == 2019) return "E"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2230) return "E"  ;
    if (arc_index == 2279) return "W"  ;
    if (arc_index == 2440) return "E"  ;
    if (arc_index == 2459) return "H"  ;
    if (arc_index == 2540) return "W"  ;
    if (arc_index == 2614) return "H"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2747) return "H"  ;
    if (arc_index == 2755) return "H"  ;
    if (arc_index == 2842) return "H"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 8)) begin 
    if (arc_index == 30) return "H"  ;
    if (arc_index == 64) return "H"  ;
    if (arc_index == 161) return "H"  ;
    if (arc_index == 164) return "H"  ;
    if (arc_index == 175) return "H"  ;
    if (arc_index == 177) return "H"  ;
    if (arc_index == 199) return "H"  ;
    if (arc_index == 203) return "E"  ;
    if (arc_index == 208) return "E"  ;
    if (arc_index == 213) return "E"  ;
    if (arc_index == 215) return "E"  ;
    if (arc_index == 220) return "E"  ;
    if (arc_index == 228) return "W"  ;
    if (arc_index == 231) return "W"  ;
    if (arc_index == 242) return "W"  ;
    if (arc_index == 244) return "W"  ;
    if (arc_index == 245) return "H"  ;
    if (arc_index == 249) return "H"  ;
    if (arc_index == 250) return "H"  ;
    if (arc_index == 252) return "H"  ;
    if (arc_index == 253) return "H"  ;
    if (arc_index == 255) return "H"  ;
    if (arc_index == 257) return "H"  ;
    if (arc_index == 260) return "H"  ;
    if (arc_index == 261) return "W"  ;
    if (arc_index == 275) return "W"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 311) return "W"  ;
    if (arc_index == 312) return "W"  ;
    if (arc_index == 315) return "W"  ;
    if (arc_index == 320) return "W"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 323) return "W"  ;
    if (arc_index == 325) return "W"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 329) return "W"  ;
    if (arc_index == 354) return "E"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 420) return "H"  ;
    if (arc_index == 442) return "H"  ;
    if (arc_index == 528) return "H"  ;
    if (arc_index == 552) return "E"  ;
    if (arc_index == 556) return "E"  ;
    if (arc_index == 566) return "E"  ;
    if (arc_index == 568) return "E"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 617) return "H"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 634) return "W"  ;
    if (arc_index == 649) return "E"  ;
    if (arc_index == 660) return "H"  ;
    if (arc_index == 682) return "E"  ;
    if (arc_index == 683) return "E"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 685) return "W"  ;
    if (arc_index == 686) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 688) return "W"  ;
    if (arc_index == 689) return "W"  ;
    if (arc_index == 690) return "W"  ;
    if (arc_index == 691) return "W"  ;
    if (arc_index == 692) return "W"  ;
    if (arc_index == 693) return "W"  ;
    if (arc_index == 694) return "E"  ;
    if (arc_index == 695) return "E"  ;
    if (arc_index == 696) return "E"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 698) return "W"  ;
    if (arc_index == 699) return "W"  ;
    if (arc_index == 700) return "W"  ;
    if (arc_index == 701) return "W"  ;
    if (arc_index == 702) return "W"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 710) return "W"  ;
    if (arc_index == 715) return "H"  ;
    if (arc_index == 721) return "H"  ;
    if (arc_index == 760) return "H"  ;
    if (arc_index == 762) return "E"  ;
    if (arc_index == 814) return "W"  ;
    if (arc_index == 827) return "W"  ;
    if (arc_index == 842) return "E"  ;
    if (arc_index == 846) return "E"  ;
    if (arc_index == 847) return "E"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 959) return "H"  ;
    if (arc_index == 1016) return "H"  ;
    if (arc_index == 1118) return "H"  ;
    if (arc_index == 1136) return "H"  ;
    if (arc_index == 1174) return "E"  ;
    if (arc_index == 1220) return "H"  ;
    if (arc_index == 1239) return "H"  ;
    if (arc_index == 1251) return "H"  ;
    if (arc_index == 1259) return "H"  ;
    if (arc_index == 1263) return "E"  ;
    if (arc_index == 1329) return "H"  ;
    if (arc_index == 1379) return "E"  ;
    if (arc_index == 1409) return "E"  ;
    if (arc_index == 1414) return "E"  ;
    if (arc_index == 1420) return "E"  ;
    if (arc_index == 1426) return "E"  ;
    if (arc_index == 1445) return "H"  ;
    if (arc_index == 1458) return "E"  ;
    if (arc_index == 1501) return "E"  ;
    if (arc_index == 1534) return "H"  ;
    if (arc_index == 1548) return "H"  ;
    if (arc_index == 1558) return "W"  ;
    if (arc_index == 1583) return "W"  ;
    if (arc_index == 1653) return "W"  ;
    if (arc_index == 1679) return "H"  ;
    if (arc_index == 1685) return "H"  ;
    if (arc_index == 1688) return "W"  ;
    if (arc_index == 1705) return "W"  ;
    if (arc_index == 1708) return "W"  ;
    if (arc_index == 1714) return "E"  ;
    if (arc_index == 1763) return "E"  ;
    if (arc_index == 1775) return "E"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1778) return "W"  ;
    if (arc_index == 1793) return "W"  ;
    if (arc_index == 1825) return "E"  ;
    if (arc_index == 1832) return "H"  ;
    if (arc_index == 1895) return "E"  ;
    if (arc_index == 1978) return "E"  ;
    if (arc_index == 2068) return "E"  ;
    if (arc_index == 2090) return "E"  ;
    if (arc_index == 2091) return "E"  ;
    if (arc_index == 2093) return "W"  ;
    if (arc_index == 2095) return "W"  ;
    if (arc_index == 2097) return "W"  ;
    if (arc_index == 2098) return "W"  ;
    if (arc_index == 2100) return "W"  ;
    if (arc_index == 2103) return "W"  ;
    if (arc_index == 2104) return "W"  ;
    if (arc_index == 2106) return "W"  ;
    if (arc_index == 2108) return "W"  ;
    if (arc_index == 2123) return "W"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2196) return "W"  ;
    if (arc_index == 2214) return "W"  ;
    if (arc_index == 2262) return "E"  ;
    if (arc_index == 2295) return "E"  ;
    if (arc_index == 2329) return "E"  ;
    if (arc_index == 2335) return "W"  ;
    if (arc_index == 2340) return "W"  ;
    if (arc_index == 2341) return "W"  ;
    if (arc_index == 2342) return "W"  ;
    if (arc_index == 2346) return "W"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2367) return "W"  ;
    if (arc_index == 2380) return "W"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2424) return "W"  ;
    if (arc_index == 2467) return "E"  ;
    if (arc_index == 2471) return "E"  ;
    if (arc_index == 2481) return "H"  ;
    if (arc_index == 2490) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2601) return "E"  ;
    if (arc_index == 2605) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2635) return "W"  ;
    if (arc_index == 2636) return "H"  ;
    if (arc_index == 2637) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2757) return "E"  ;
    if (arc_index == 2769) return "H"  ;
    if (arc_index == 2777) return "H"  ;
    if (arc_index == 2786) return "E"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2864) return "H"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2906) return "E"  ;
    if (arc_index == 2916) return "E"  ;
    if (arc_index == 2923) return "W"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 10)) begin 
    if (arc_index == 86) return "H"  ;
    if (arc_index == 197) return "H"  ;
    if (arc_index == 254) return "H"  ;
    if (arc_index == 267) return "H"  ;
    if (arc_index == 314) return "H"  ;
    if (arc_index == 442) return "H"  ;
    if (arc_index == 563) return "H"  ;
    if (arc_index == 621) return "W"  ;
    if (arc_index == 628) return "W"  ;
    if (arc_index == 639) return "H"  ;
    if (arc_index == 682) return "H"  ;
    if (arc_index == 704) return "H"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 707) return "W"  ;
    if (arc_index == 708) return "W"  ;
    if (arc_index == 709) return "W"  ;
    if (arc_index == 710) return "W"  ;
    if (arc_index == 711) return "W"  ;
    if (arc_index == 712) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 714) return "W"  ;
    if (arc_index == 715) return "W"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 718) return "W"  ;
    if (arc_index == 719) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 721) return "W"  ;
    if (arc_index == 722) return "W"  ;
    if (arc_index == 723) return "W"  ;
    if (arc_index == 724) return "W"  ;
    if (arc_index == 725) return "W"  ;
    if (arc_index == 737) return "H"  ;
    if (arc_index == 782) return "H"  ;
    if (arc_index == 981) return "H"  ;
    if (arc_index == 1158) return "H"  ;
    if (arc_index == 1242) return "H"  ;
    if (arc_index == 1346) return "H"  ;
    if (arc_index == 1351) return "H"  ;
    if (arc_index == 1467) return "H"  ;
    if (arc_index == 1468) return "H"  ;
    if (arc_index == 1547) return "W"  ;
    if (arc_index == 1556) return "H"  ;
    if (arc_index == 1570) return "H"  ;
    if (arc_index == 1701) return "H"  ;
    if (arc_index == 1766) return "H"  ;
    if (arc_index == 1854) return "H"  ;
    if (arc_index == 2101) return "H"  ;
    if (arc_index == 2105) return "H"  ;
    if (arc_index == 2111) return "H"  ;
    if (arc_index == 2503) return "H"  ;
    if (arc_index == 2596) return "H"  ;
    if (arc_index == 2616) return "H"  ;
    if (arc_index == 2626) return "W"  ;
    if (arc_index == 2628) return "W"  ;
    if (arc_index == 2629) return "W"  ;
    if (arc_index == 2658) return "H"  ;
    if (arc_index == 2791) return "H"  ;
    if (arc_index == 2799) return "H"  ;
    if (arc_index == 2886) return "H"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 8)) begin 
    if (arc_index == 108) return "H"  ;
    if (arc_index == 219) return "H"  ;
    if (arc_index == 240) return "W"  ;
    if (arc_index == 252) return "E"  ;
    if (arc_index == 289) return "H"  ;
    if (arc_index == 361) return "E"  ;
    if (arc_index == 435) return "E"  ;
    if (arc_index == 464) return "H"  ;
    if (arc_index == 620) return "W"  ;
    if (arc_index == 661) return "H"  ;
    if (arc_index == 680) return "E"  ;
    if (arc_index == 704) return "H"  ;
    if (arc_index == 726) return "H"  ;
    if (arc_index == 727) return "W"  ;
    if (arc_index == 728) return "W"  ;
    if (arc_index == 729) return "W"  ;
    if (arc_index == 730) return "W"  ;
    if (arc_index == 731) return "E"  ;
    if (arc_index == 732) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 735) return "W"  ;
    if (arc_index == 736) return "W"  ;
    if (arc_index == 737) return "W"  ;
    if (arc_index == 738) return "W"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 740) return "W"  ;
    if (arc_index == 741) return "W"  ;
    if (arc_index == 742) return "W"  ;
    if (arc_index == 743) return "W"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 746) return "W"  ;
    if (arc_index == 747) return "W"  ;
    if (arc_index == 759) return "H"  ;
    if (arc_index == 804) return "H"  ;
    if (arc_index == 860) return "H"  ;
    if (arc_index == 861) return "E"  ;
    if (arc_index == 864) return "E"  ;
    if (arc_index == 867) return "E"  ;
    if (arc_index == 871) return "E"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 1003) return "H"  ;
    if (arc_index == 1043) return "W"  ;
    if (arc_index == 1135) return "W"  ;
    if (arc_index == 1180) return "H"  ;
    if (arc_index == 1248) return "W"  ;
    if (arc_index == 1264) return "H"  ;
    if (arc_index == 1307) return "W"  ;
    if (arc_index == 1342) return "W"  ;
    if (arc_index == 1369) return "W"  ;
    if (arc_index == 1373) return "H"  ;
    if (arc_index == 1489) return "H"  ;
    if (arc_index == 1497) return "E"  ;
    if (arc_index == 1513) return "E"  ;
    if (arc_index == 1562) return "E"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1565) return "W"  ;
    if (arc_index == 1568) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1574) return "W"  ;
    if (arc_index == 1578) return "H"  ;
    if (arc_index == 1592) return "H"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1723) return "H"  ;
    if (arc_index == 1876) return "H"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2016) return "E"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2209) return "E"  ;
    if (arc_index == 2428) return "E"  ;
    if (arc_index == 2525) return "H"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2646) return "W"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2657) return "W"  ;
    if (arc_index == 2660) return "W"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2680) return "H"  ;
    if (arc_index == 2813) return "H"  ;
    if (arc_index == 2821) return "H"  ;
    if (arc_index == 2908) return "H"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 4)) begin 
    if (arc_index == 4) return "H"  ;
    if (arc_index == 95) return "W"  ;
    if (arc_index == 123) return "W"  ;
    if (arc_index == 130) return "H"  ;
    if (arc_index == 189) return "H"  ;
    if (arc_index == 241) return "H"  ;
    if (arc_index == 247) return "W"  ;
    if (arc_index == 248) return "W"  ;
    if (arc_index == 256) return "W"  ;
    if (arc_index == 262) return "W"  ;
    if (arc_index == 263) return "W"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 311) return "H"  ;
    if (arc_index == 333) return "H"  ;
    if (arc_index == 340) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 384) return "W"  ;
    if (arc_index == 486) return "H"  ;
    if (arc_index == 493) return "H"  ;
    if (arc_index == 560) return "H"  ;
    if (arc_index == 570) return "H"  ;
    if (arc_index == 609) return "H"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 664) return "W"  ;
    if (arc_index == 683) return "H"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 726) return "H"  ;
    if (arc_index == 748) return "H"  ;
    if (arc_index == 749) return "E"  ;
    if (arc_index == 750) return "E"  ;
    if (arc_index == 751) return "W"  ;
    if (arc_index == 752) return "W"  ;
    if (arc_index == 753) return "W"  ;
    if (arc_index == 754) return "W"  ;
    if (arc_index == 755) return "W"  ;
    if (arc_index == 756) return "W"  ;
    if (arc_index == 757) return "W"  ;
    if (arc_index == 758) return "W"  ;
    if (arc_index == 759) return "W"  ;
    if (arc_index == 760) return "E"  ;
    if (arc_index == 761) return "E"  ;
    if (arc_index == 762) return "E"  ;
    if (arc_index == 763) return "E"  ;
    if (arc_index == 764) return "E"  ;
    if (arc_index == 765) return "E"  ;
    if (arc_index == 766) return "W"  ;
    if (arc_index == 767) return "W"  ;
    if (arc_index == 768) return "E"  ;
    if (arc_index == 769) return "E"  ;
    if (arc_index == 771) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 775) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 780) return "E"  ;
    if (arc_index == 781) return "H"  ;
    if (arc_index == 782) return "E"  ;
    if (arc_index == 784) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 826) return "H"  ;
    if (arc_index == 843) return "H"  ;
    if (arc_index == 889) return "E"  ;
    if (arc_index == 949) return "E"  ;
    if (arc_index == 950) return "E"  ;
    if (arc_index == 996) return "E"  ;
    if (arc_index == 1025) return "H"  ;
    if (arc_index == 1047) return "H"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1062) return "W"  ;
    if (arc_index == 1120) return "W"  ;
    if (arc_index == 1197) return "W"  ;
    if (arc_index == 1202) return "H"  ;
    if (arc_index == 1286) return "H"  ;
    if (arc_index == 1388) return "H"  ;
    if (arc_index == 1389) return "W"  ;
    if (arc_index == 1391) return "W"  ;
    if (arc_index == 1395) return "H"  ;
    if (arc_index == 1400) return "W"  ;
    if (arc_index == 1406) return "W"  ;
    if (arc_index == 1424) return "W"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1454) return "W"  ;
    if (arc_index == 1459) return "W"  ;
    if (arc_index == 1476) return "W"  ;
    if (arc_index == 1511) return "H"  ;
    if (arc_index == 1600) return "H"  ;
    if (arc_index == 1614) return "H"  ;
    if (arc_index == 1629) return "H"  ;
    if (arc_index == 1645) return "H"  ;
    if (arc_index == 1663) return "E"  ;
    if (arc_index == 1709) return "W"  ;
    if (arc_index == 1715) return "W"  ;
    if (arc_index == 1727) return "W"  ;
    if (arc_index == 1738) return "E"  ;
    if (arc_index == 1745) return "H"  ;
    if (arc_index == 1751) return "H"  ;
    if (arc_index == 1755) return "H"  ;
    if (arc_index == 1757) return "E"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1762) return "W"  ;
    if (arc_index == 1771) return "W"  ;
    if (arc_index == 1800) return "W"  ;
    if (arc_index == 1816) return "W"  ;
    if (arc_index == 1838) return "E"  ;
    if (arc_index == 1840) return "E"  ;
    if (arc_index == 1866) return "E"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1898) return "H"  ;
    if (arc_index == 1933) return "H"  ;
    if (arc_index == 1946) return "H"  ;
    if (arc_index == 1999) return "H"  ;
    if (arc_index == 2025) return "E"  ;
    if (arc_index == 2026) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2033) return "E"  ;
    if (arc_index == 2041) return "E"  ;
    if (arc_index == 2057) return "W"  ;
    if (arc_index == 2102) return "W"  ;
    if (arc_index == 2148) return "W"  ;
    if (arc_index == 2149) return "E"  ;
    if (arc_index == 2154) return "E"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2290) return "W"  ;
    if (arc_index == 2291) return "W"  ;
    if (arc_index == 2297) return "W"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2301) return "W"  ;
    if (arc_index == 2305) return "W"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2457) return "W"  ;
    if (arc_index == 2487) return "W"  ;
    if (arc_index == 2501) return "W"  ;
    if (arc_index == 2510) return "W"  ;
    if (arc_index == 2547) return "H"  ;
    if (arc_index == 2554) return "H"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2564) return "E"  ;
    if (arc_index == 2565) return "E"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2604) return "W"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2691) return "E"  ;
    if (arc_index == 2702) return "H"  ;
    if (arc_index == 2707) return "H"  ;
    if (arc_index == 2724) return "H"  ;
    if (arc_index == 2728) return "H"  ;
    if (arc_index == 2731) return "E"  ;
    if (arc_index == 2732) return "E"  ;
    if (arc_index == 2736) return "E"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2742) return "E"  ;
    if (arc_index == 2744) return "E"  ;
    if (arc_index == 2749) return "E"  ;
    if (arc_index == 2750) return "E"  ;
    if (arc_index == 2774) return "E"  ;
    if (arc_index == 2778) return "E"  ;
    if (arc_index == 2780) return "W"  ;
    if (arc_index == 2781) return "W"  ;
    if (arc_index == 2782) return "E"  ;
    if (arc_index == 2783) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2785) return "E"  ;
    if (arc_index == 2787) return "W"  ;
    if (arc_index == 2788) return "W"  ;
    if (arc_index == 2789) return "W"  ;
    if (arc_index == 2793) return "W"  ;
    if (arc_index == 2805) return "W"  ;
    if (arc_index == 2816) return "W"  ;
    if (arc_index == 2835) return "H"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2841) return "E"  ;
    if (arc_index == 2843) return "H"  ;
    if (arc_index == 2845) return "H"  ;
    if (arc_index == 2846) return "H"  ;
    if (arc_index == 2847) return "H"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2849) return "E"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2855) return "E"  ;
    if (arc_index == 2864) return "E"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2873) return "E"  ;
    if (arc_index == 2890) return "W"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 2)) begin 
    if (arc_index == 26) return "H"  ;
    if (arc_index == 80) return "W"  ;
    if (arc_index == 152) return "H"  ;
    if (arc_index == 164) return "W"  ;
    if (arc_index == 263) return "H"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 333) return "H"  ;
    if (arc_index == 508) return "H"  ;
    if (arc_index == 565) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 705) return "H"  ;
    if (arc_index == 748) return "H"  ;
    if (arc_index == 770) return "H"  ;
    if (arc_index == 771) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 773) return "W"  ;
    if (arc_index == 774) return "W"  ;
    if (arc_index == 775) return "E"  ;
    if (arc_index == 776) return "W"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 778) return "E"  ;
    if (arc_index == 779) return "E"  ;
    if (arc_index == 780) return "E"  ;
    if (arc_index == 781) return "E"  ;
    if (arc_index == 782) return "E"  ;
    if (arc_index == 783) return "E"  ;
    if (arc_index == 784) return "E"  ;
    if (arc_index == 785) return "E"  ;
    if (arc_index == 786) return "W"  ;
    if (arc_index == 787) return "W"  ;
    if (arc_index == 788) return "E"  ;
    if (arc_index == 789) return "E"  ;
    if (arc_index == 790) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 803) return "H"  ;
    if (arc_index == 848) return "H"  ;
    if (arc_index == 1047) return "H"  ;
    if (arc_index == 1224) return "H"  ;
    if (arc_index == 1308) return "H"  ;
    if (arc_index == 1417) return "H"  ;
    if (arc_index == 1418) return "H"  ;
    if (arc_index == 1425) return "W"  ;
    if (arc_index == 1533) return "H"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1622) return "H"  ;
    if (arc_index == 1636) return "H"  ;
    if (arc_index == 1713) return "W"  ;
    if (arc_index == 1721) return "W"  ;
    if (arc_index == 1767) return "H"  ;
    if (arc_index == 1920) return "H"  ;
    if (arc_index == 2045) return "W"  ;
    if (arc_index == 2110) return "W"  ;
    if (arc_index == 2232) return "E"  ;
    if (arc_index == 2290) return "W"  ;
    if (arc_index == 2487) return "W"  ;
    if (arc_index == 2530) return "W"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2554) return "E"  ;
    if (arc_index == 2558) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2560) return "E"  ;
    if (arc_index == 2562) return "E"  ;
    if (arc_index == 2563) return "E"  ;
    if (arc_index == 2564) return "E"  ;
    if (arc_index == 2565) return "E"  ;
    if (arc_index == 2568) return "E"  ;
    if (arc_index == 2569) return "H"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2724) return "H"  ;
    if (arc_index == 2737) return "E"  ;
    if (arc_index == 2829) return "W"  ;
    if (arc_index == 2838) return "W"  ;
    if (arc_index == 2851) return "W"  ;
    if (arc_index == 2857) return "H"  ;
    if (arc_index == 2859) return "W"  ;
    if (arc_index == 2865) return "H"  ;
    if (arc_index == 2871) return "E"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 2)) begin 
    if (arc_index == 48) return "H"  ;
    if (arc_index == 73) return "H"  ;
    if (arc_index == 102) return "W"  ;
    if (arc_index == 144) return "W"  ;
    if (arc_index == 174) return "H"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 285) return "H"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 355) return "H"  ;
    if (arc_index == 411) return "W"  ;
    if (arc_index == 417) return "W"  ;
    if (arc_index == 418) return "W"  ;
    if (arc_index == 513) return "E"  ;
    if (arc_index == 530) return "H"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 645) return "W"  ;
    if (arc_index == 662) return "W"  ;
    if (arc_index == 681) return "W"  ;
    if (arc_index == 727) return "H"  ;
    if (arc_index == 770) return "H"  ;
    if (arc_index == 792) return "H"  ;
    if (arc_index == 793) return "E"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 795) return "E"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 797) return "E"  ;
    if (arc_index == 798) return "W"  ;
    if (arc_index == 799) return "W"  ;
    if (arc_index == 800) return "W"  ;
    if (arc_index == 801) return "W"  ;
    if (arc_index == 802) return "W"  ;
    if (arc_index == 803) return "W"  ;
    if (arc_index == 804) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 806) return "E"  ;
    if (arc_index == 807) return "E"  ;
    if (arc_index == 808) return "E"  ;
    if (arc_index == 809) return "E"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 811) return "E"  ;
    if (arc_index == 812) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 825) return "H"  ;
    if (arc_index == 859) return "H"  ;
    if (arc_index == 870) return "H"  ;
    if (arc_index == 925) return "E"  ;
    if (arc_index == 927) return "E"  ;
    if (arc_index == 934) return "E"  ;
    if (arc_index == 936) return "E"  ;
    if (arc_index == 1011) return "E"  ;
    if (arc_index == 1069) return "H"  ;
    if (arc_index == 1123) return "H"  ;
    if (arc_index == 1246) return "H"  ;
    if (arc_index == 1330) return "H"  ;
    if (arc_index == 1372) return "H"  ;
    if (arc_index == 1439) return "H"  ;
    if (arc_index == 1447) return "W"  ;
    if (arc_index == 1528) return "E"  ;
    if (arc_index == 1555) return "H"  ;
    if (arc_index == 1644) return "H"  ;
    if (arc_index == 1658) return "H"  ;
    if (arc_index == 1740) return "H"  ;
    if (arc_index == 1789) return "H"  ;
    if (arc_index == 1937) return "H"  ;
    if (arc_index == 1942) return "H"  ;
    if (arc_index == 2002) return "H"  ;
    if (arc_index == 2004) return "H"  ;
    if (arc_index == 2006) return "H"  ;
    if (arc_index == 2007) return "H"  ;
    if (arc_index == 2012) return "H"  ;
    if (arc_index == 2013) return "H"  ;
    if (arc_index == 2014) return "H"  ;
    if (arc_index == 2015) return "H"  ;
    if (arc_index == 2020) return "H"  ;
    if (arc_index == 2021) return "H"  ;
    if (arc_index == 2023) return "H"  ;
    if (arc_index == 2035) return "H"  ;
    if (arc_index == 2067) return "W"  ;
    if (arc_index == 2137) return "W"  ;
    if (arc_index == 2230) return "W"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2456) return "W"  ;
    if (arc_index == 2509) return "W"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2577) return "E"  ;
    if (arc_index == 2578) return "E"  ;
    if (arc_index == 2584) return "E"  ;
    if (arc_index == 2586) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2588) return "E"  ;
    if (arc_index == 2591) return "H"  ;
    if (arc_index == 2592) return "E"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2746) return "H"  ;
    if (arc_index == 2747) return "E"  ;
    if (arc_index == 2765) return "E"  ;
    if (arc_index == 2854) return "E"  ;
    if (arc_index == 2868) return "E"  ;
    if (arc_index == 2879) return "H"  ;
    if (arc_index == 2887) return "H"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 9)) begin 
    if (arc_index == 11) return "E"  ;
    if (arc_index == 53) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 70) return "H"  ;
    if (arc_index == 109) return "H"  ;
    if (arc_index == 124) return "H"  ;
    if (arc_index == 169) return "H"  ;
    if (arc_index == 196) return "H"  ;
    if (arc_index == 203) return "H"  ;
    if (arc_index == 215) return "E"  ;
    if (arc_index == 255) return "E"  ;
    if (arc_index == 267) return "E"  ;
    if (arc_index == 272) return "E"  ;
    if (arc_index == 301) return "W"  ;
    if (arc_index == 307) return "H"  ;
    if (arc_index == 308) return "H"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 326) return "W"  ;
    if (arc_index == 327) return "W"  ;
    if (arc_index == 377) return "H"  ;
    if (arc_index == 432) return "E"  ;
    if (arc_index == 433) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 536) return "E"  ;
    if (arc_index == 552) return "H"  ;
    if (arc_index == 566) return "H"  ;
    if (arc_index == 568) return "E"  ;
    if (arc_index == 601) return "W"  ;
    if (arc_index == 619) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 635) return "W"  ;
    if (arc_index == 667) return "W"  ;
    if (arc_index == 685) return "W"  ;
    if (arc_index == 701) return "W"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 749) return "H"  ;
    if (arc_index == 792) return "H"  ;
    if (arc_index == 814) return "W"  ;
    if (arc_index == 815) return "W"  ;
    if (arc_index == 816) return "W"  ;
    if (arc_index == 817) return "W"  ;
    if (arc_index == 818) return "W"  ;
    if (arc_index == 819) return "W"  ;
    if (arc_index == 820) return "W"  ;
    if (arc_index == 821) return "W"  ;
    if (arc_index == 822) return "W"  ;
    if (arc_index == 823) return "W"  ;
    if (arc_index == 824) return "E"  ;
    if (arc_index == 825) return "E"  ;
    if (arc_index == 826) return "W"  ;
    if (arc_index == 827) return "W"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 830) return "E"  ;
    if (arc_index == 831) return "W"  ;
    if (arc_index == 832) return "W"  ;
    if (arc_index == 833) return "W"  ;
    if (arc_index == 834) return "W"  ;
    if (arc_index == 835) return "E"  ;
    if (arc_index == 842) return "E"  ;
    if (arc_index == 844) return "E"  ;
    if (arc_index == 847) return "H"  ;
    if (arc_index == 892) return "H"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 1037) return "W"  ;
    if (arc_index == 1070) return "W"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1091) return "H"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1142) return "W"  ;
    if (arc_index == 1146) return "W"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1205) return "W"  ;
    if (arc_index == 1253) return "W"  ;
    if (arc_index == 1268) return "H"  ;
    if (arc_index == 1316) return "W"  ;
    if (arc_index == 1323) return "W"  ;
    if (arc_index == 1343) return "W"  ;
    if (arc_index == 1344) return "W"  ;
    if (arc_index == 1345) return "W"  ;
    if (arc_index == 1348) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1352) return "H"  ;
    if (arc_index == 1353) return "H"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1359) return "W"  ;
    if (arc_index == 1362) return "W"  ;
    if (arc_index == 1363) return "W"  ;
    if (arc_index == 1375) return "E"  ;
    if (arc_index == 1404) return "E"  ;
    if (arc_index == 1420) return "E"  ;
    if (arc_index == 1421) return "E"  ;
    if (arc_index == 1461) return "H"  ;
    if (arc_index == 1482) return "E"  ;
    if (arc_index == 1491) return "E"  ;
    if (arc_index == 1493) return "E"  ;
    if (arc_index == 1552) return "W"  ;
    if (arc_index == 1558) return "W"  ;
    if (arc_index == 1577) return "H"  ;
    if (arc_index == 1583) return "W"  ;
    if (arc_index == 1588) return "W"  ;
    if (arc_index == 1613) return "W"  ;
    if (arc_index == 1619) return "E"  ;
    if (arc_index == 1666) return "H"  ;
    if (arc_index == 1680) return "H"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1769) return "E"  ;
    if (arc_index == 1770) return "E"  ;
    if (arc_index == 1774) return "E"  ;
    if (arc_index == 1780) return "E"  ;
    if (arc_index == 1796) return "E"  ;
    if (arc_index == 1811) return "H"  ;
    if (arc_index == 1852) return "H"  ;
    if (arc_index == 1880) return "E"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1964) return "H"  ;
    if (arc_index == 1989) return "E"  ;
    if (arc_index == 1996) return "E"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2068) return "E"  ;
    if (arc_index == 2070) return "E"  ;
    if (arc_index == 2089) return "E"  ;
    if (arc_index == 2092) return "E"  ;
    if (arc_index == 2100) return "E"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2192) return "E"  ;
    if (arc_index == 2196) return "E"  ;
    if (arc_index == 2198) return "W"  ;
    if (arc_index == 2267) return "W"  ;
    if (arc_index == 2286) return "E"  ;
    if (arc_index == 2289) return "E"  ;
    if (arc_index == 2295) return "E"  ;
    if (arc_index == 2310) return "E"  ;
    if (arc_index == 2326) return "W"  ;
    if (arc_index == 2332) return "W"  ;
    if (arc_index == 2333) return "W"  ;
    if (arc_index == 2336) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2343) return "W"  ;
    if (arc_index == 2344) return "W"  ;
    if (arc_index == 2345) return "W"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2351) return "W"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2365) return "W"  ;
    if (arc_index == 2379) return "W"  ;
    if (arc_index == 2407) return "W"  ;
    if (arc_index == 2410) return "W"  ;
    if (arc_index == 2467) return "E"  ;
    if (arc_index == 2492) return "E"  ;
    if (arc_index == 2599) return "E"  ;
    if (arc_index == 2600) return "W"  ;
    if (arc_index == 2606) return "W"  ;
    if (arc_index == 2611) return "W"  ;
    if (arc_index == 2613) return "H"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2615) return "W"  ;
    if (arc_index == 2624) return "W"  ;
    if (arc_index == 2634) return "W"  ;
    if (arc_index == 2703) return "W"  ;
    if (arc_index == 2768) return "H"  ;
    if (arc_index == 2775) return "H"  ;
    if (arc_index == 2776) return "H"  ;
    if (arc_index == 2830) return "H"  ;
    if (arc_index == 2833) return "E"  ;
    if (arc_index == 2836) return "E"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2882) return "E"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2901) return "H"  ;
    if (arc_index == 2904) return "H"  ;
    if (arc_index == 2909) return "H"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2912) return "W"  ;
    if (arc_index == 2915) return "W"  ;
    if (arc_index == 2918) return "W"  ;
    if (arc_index == 2919) return "W"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 6)) begin 
    if (arc_index == 4) return "W"  ;
    if (arc_index == 5) return "H"  ;
    if (arc_index == 9) return "E"  ;
    if (arc_index == 92) return "H"  ;
    if (arc_index == 95) return "H"  ;
    if (arc_index == 113) return "H"  ;
    if (arc_index == 125) return "E"  ;
    if (arc_index == 200) return "W"  ;
    if (arc_index == 202) return "W"  ;
    if (arc_index == 204) return "W"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 207) return "W"  ;
    if (arc_index == 211) return "W"  ;
    if (arc_index == 212) return "W"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 218) return "H"  ;
    if (arc_index == 244) return "W"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 311) return "W"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 323) return "W"  ;
    if (arc_index == 325) return "W"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 329) return "H"  ;
    if (arc_index == 340) return "H"  ;
    if (arc_index == 399) return "H"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 436) return "E"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 475) return "E"  ;
    if (arc_index == 480) return "E"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 512) return "E"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 547) return "W"  ;
    if (arc_index == 553) return "W"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 574) return "H"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 601) return "W"  ;
    if (arc_index == 613) return "W"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 642) return "W"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 688) return "W"  ;
    if (arc_index == 690) return "W"  ;
    if (arc_index == 691) return "W"  ;
    if (arc_index == 693) return "W"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 698) return "W"  ;
    if (arc_index == 699) return "W"  ;
    if (arc_index == 758) return "E"  ;
    if (arc_index == 760) return "E"  ;
    if (arc_index == 762) return "E"  ;
    if (arc_index == 771) return "H"  ;
    if (arc_index == 772) return "H"  ;
    if (arc_index == 791) return "H"  ;
    if (arc_index == 814) return "H"  ;
    if (arc_index == 826) return "W"  ;
    if (arc_index == 836) return "W"  ;
    if (arc_index == 837) return "W"  ;
    if (arc_index == 838) return "W"  ;
    if (arc_index == 839) return "W"  ;
    if (arc_index == 840) return "W"  ;
    if (arc_index == 841) return "E"  ;
    if (arc_index == 842) return "E"  ;
    if (arc_index == 843) return "E"  ;
    if (arc_index == 844) return "E"  ;
    if (arc_index == 845) return "E"  ;
    if (arc_index == 846) return "E"  ;
    if (arc_index == 847) return "E"  ;
    if (arc_index == 848) return "W"  ;
    if (arc_index == 849) return "W"  ;
    if (arc_index == 850) return "W"  ;
    if (arc_index == 851) return "W"  ;
    if (arc_index == 852) return "W"  ;
    if (arc_index == 853) return "W"  ;
    if (arc_index == 854) return "W"  ;
    if (arc_index == 855) return "W"  ;
    if (arc_index == 856) return "E"  ;
    if (arc_index == 857) return "E"  ;
    if (arc_index == 863) return "E"  ;
    if (arc_index == 869) return "H"  ;
    if (arc_index == 892) return "E"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 901) return "E"  ;
    if (arc_index == 914) return "H"  ;
    if (arc_index == 945) return "H"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 961) return "E"  ;
    if (arc_index == 971) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1076) return "W"  ;
    if (arc_index == 1094) return "W"  ;
    if (arc_index == 1113) return "H"  ;
    if (arc_index == 1120) return "H"  ;
    if (arc_index == 1124) return "W"  ;
    if (arc_index == 1174) return "E"  ;
    if (arc_index == 1190) return "E"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1286) return "E"  ;
    if (arc_index == 1290) return "H"  ;
    if (arc_index == 1321) return "W"  ;
    if (arc_index == 1334) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1374) return "H"  ;
    if (arc_index == 1394) return "H"  ;
    if (arc_index == 1399) return "E"  ;
    if (arc_index == 1401) return "E"  ;
    if (arc_index == 1404) return "E"  ;
    if (arc_index == 1405) return "E"  ;
    if (arc_index == 1410) return "E"  ;
    if (arc_index == 1411) return "W"  ;
    if (arc_index == 1413) return "W"  ;
    if (arc_index == 1414) return "E"  ;
    if (arc_index == 1415) return "E"  ;
    if (arc_index == 1421) return "E"  ;
    if (arc_index == 1422) return "E"  ;
    if (arc_index == 1423) return "E"  ;
    if (arc_index == 1427) return "E"  ;
    if (arc_index == 1428) return "W"  ;
    if (arc_index == 1430) return "W"  ;
    if (arc_index == 1452) return "W"  ;
    if (arc_index == 1455) return "W"  ;
    if (arc_index == 1456) return "W"  ;
    if (arc_index == 1460) return "E"  ;
    if (arc_index == 1461) return "E"  ;
    if (arc_index == 1462) return "E"  ;
    if (arc_index == 1470) return "E"  ;
    if (arc_index == 1471) return "E"  ;
    if (arc_index == 1476) return "W"  ;
    if (arc_index == 1483) return "H"  ;
    if (arc_index == 1485) return "H"  ;
    if (arc_index == 1492) return "W"  ;
    if (arc_index == 1498) return "W"  ;
    if (arc_index == 1530) return "W"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1543) return "W"  ;
    if (arc_index == 1558) return "W"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1599) return "H"  ;
    if (arc_index == 1624) return "E"  ;
    if (arc_index == 1670) return "E"  ;
    if (arc_index == 1688) return "H"  ;
    if (arc_index == 1702) return "H"  ;
    if (arc_index == 1704) return "H"  ;
    if (arc_index == 1729) return "H"  ;
    if (arc_index == 1739) return "E"  ;
    if (arc_index == 1760) return "E"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1773) return "W"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1793) return "E"  ;
    if (arc_index == 1800) return "E"  ;
    if (arc_index == 1816) return "E"  ;
    if (arc_index == 1828) return "E"  ;
    if (arc_index == 1833) return "H"  ;
    if (arc_index == 1862) return "H"  ;
    if (arc_index == 1895) return "E"  ;
    if (arc_index == 1906) return "E"  ;
    if (arc_index == 1959) return "W"  ;
    if (arc_index == 1971) return "W"  ;
    if (arc_index == 1985) return "W"  ;
    if (arc_index == 1986) return "H"  ;
    if (arc_index == 1997) return "E"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2055) return "E"  ;
    if (arc_index == 2093) return "W"  ;
    if (arc_index == 2097) return "W"  ;
    if (arc_index == 2104) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2152) return "E"  ;
    if (arc_index == 2171) return "E"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2215) return "W"  ;
    if (arc_index == 2252) return "W"  ;
    if (arc_index == 2260) return "W"  ;
    if (arc_index == 2262) return "E"  ;
    if (arc_index == 2265) return "W"  ;
    if (arc_index == 2268) return "W"  ;
    if (arc_index == 2274) return "W"  ;
    if (arc_index == 2302) return "W"  ;
    if (arc_index == 2318) return "W"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2449) return "W"  ;
    if (arc_index == 2467) return "E"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2471) return "E"  ;
    if (arc_index == 2476) return "E"  ;
    if (arc_index == 2481) return "E"  ;
    if (arc_index == 2482) return "E"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2504) return "E"  ;
    if (arc_index == 2506) return "E"  ;
    if (arc_index == 2531) return "E"  ;
    if (arc_index == 2538) return "E"  ;
    if (arc_index == 2543) return "E"  ;
    if (arc_index == 2548) return "E"  ;
    if (arc_index == 2550) return "E"  ;
    if (arc_index == 2554) return "E"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2603) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2608) return "W"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2635) return "H"  ;
    if (arc_index == 2687) return "E"  ;
    if (arc_index == 2757) return "E"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2779) return "E"  ;
    if (arc_index == 2782) return "E"  ;
    if (arc_index == 2786) return "E"  ;
    if (arc_index == 2790) return "H"  ;
    if (arc_index == 2794) return "H"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2832) return "W"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2862) return "E"  ;
    if (arc_index == 2923) return "H"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 6)) begin 
    if (arc_index == 19) return "H"  ;
    if (arc_index == 27) return "H"  ;
    if (arc_index == 114) return "H"  ;
    if (arc_index == 139) return "E"  ;
    if (arc_index == 146) return "E"  ;
    if (arc_index == 147) return "E"  ;
    if (arc_index == 150) return "E"  ;
    if (arc_index == 240) return "H"  ;
    if (arc_index == 351) return "H"  ;
    if (arc_index == 392) return "E"  ;
    if (arc_index == 396) return "E"  ;
    if (arc_index == 416) return "E"  ;
    if (arc_index == 421) return "H"  ;
    if (arc_index == 429) return "W"  ;
    if (arc_index == 595) return "W"  ;
    if (arc_index == 596) return "H"  ;
    if (arc_index == 661) return "E"  ;
    if (arc_index == 671) return "E"  ;
    if (arc_index == 680) return "E"  ;
    if (arc_index == 727) return "W"  ;
    if (arc_index == 728) return "W"  ;
    if (arc_index == 732) return "W"  ;
    if (arc_index == 738) return "W"  ;
    if (arc_index == 793) return "H"  ;
    if (arc_index == 804) return "E"  ;
    if (arc_index == 836) return "H"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 859) return "W"  ;
    if (arc_index == 860) return "E"  ;
    if (arc_index == 861) return "E"  ;
    if (arc_index == 862) return "E"  ;
    if (arc_index == 863) return "E"  ;
    if (arc_index == 864) return "E"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 866) return "W"  ;
    if (arc_index == 867) return "E"  ;
    if (arc_index == 868) return "E"  ;
    if (arc_index == 869) return "E"  ;
    if (arc_index == 870) return "W"  ;
    if (arc_index == 871) return "E"  ;
    if (arc_index == 872) return "E"  ;
    if (arc_index == 873) return "E"  ;
    if (arc_index == 874) return "E"  ;
    if (arc_index == 875) return "W"  ;
    if (arc_index == 876) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 878) return "W"  ;
    if (arc_index == 879) return "W"  ;
    if (arc_index == 891) return "H"  ;
    if (arc_index == 927) return "E"  ;
    if (arc_index == 936) return "H"  ;
    if (arc_index == 1043) return "W"  ;
    if (arc_index == 1114) return "W"  ;
    if (arc_index == 1129) return "W"  ;
    if (arc_index == 1135) return "H"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1248) return "W"  ;
    if (arc_index == 1258) return "W"  ;
    if (arc_index == 1307) return "W"  ;
    if (arc_index == 1312) return "H"  ;
    if (arc_index == 1371) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1378) return "W"  ;
    if (arc_index == 1381) return "W"  ;
    if (arc_index == 1384) return "W"  ;
    if (arc_index == 1396) return "H"  ;
    if (arc_index == 1505) return "H"  ;
    if (arc_index == 1513) return "E"  ;
    if (arc_index == 1564) return "E"  ;
    if (arc_index == 1565) return "W"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1621) return "H"  ;
    if (arc_index == 1710) return "H"  ;
    if (arc_index == 1724) return "H"  ;
    if (arc_index == 1855) return "H"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2008) return "H"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2011) return "E"  ;
    if (arc_index == 2016) return "E"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2086) return "W"  ;
    if (arc_index == 2195) return "W"  ;
    if (arc_index == 2219) return "W"  ;
    if (arc_index == 2230) return "E"  ;
    if (arc_index == 2314) return "W"  ;
    if (arc_index == 2514) return "E"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2657) return "H"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2812) return "H"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 2)) begin 
    if (arc_index == 12) return "H"  ;
    if (arc_index == 41) return "H"  ;
    if (arc_index == 49) return "H"  ;
    if (arc_index == 80) return "H"  ;
    if (arc_index == 136) return "H"  ;
    if (arc_index == 152) return "H"  ;
    if (arc_index == 211) return "H"  ;
    if (arc_index == 244) return "H"  ;
    if (arc_index == 247) return "H"  ;
    if (arc_index == 262) return "H"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 373) return "H"  ;
    if (arc_index == 443) return "H"  ;
    if (arc_index == 450) return "E"  ;
    if (arc_index == 486) return "E"  ;
    if (arc_index == 508) return "E"  ;
    if (arc_index == 550) return "E"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 618) return "H"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 751) return "W"  ;
    if (arc_index == 753) return "W"  ;
    if (arc_index == 770) return "W"  ;
    if (arc_index == 774) return "W"  ;
    if (arc_index == 779) return "W"  ;
    if (arc_index == 783) return "W"  ;
    if (arc_index == 787) return "W"  ;
    if (arc_index == 789) return "W"  ;
    if (arc_index == 803) return "W"  ;
    if (arc_index == 815) return "H"  ;
    if (arc_index == 840) return "H"  ;
    if (arc_index == 849) return "W"  ;
    if (arc_index == 858) return "H"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 880) return "W"  ;
    if (arc_index == 881) return "W"  ;
    if (arc_index == 882) return "W"  ;
    if (arc_index == 883) return "E"  ;
    if (arc_index == 884) return "E"  ;
    if (arc_index == 885) return "E"  ;
    if (arc_index == 886) return "E"  ;
    if (arc_index == 887) return "E"  ;
    if (arc_index == 888) return "E"  ;
    if (arc_index == 889) return "E"  ;
    if (arc_index == 890) return "E"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 892) return "E"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 894) return "E"  ;
    if (arc_index == 895) return "E"  ;
    if (arc_index == 896) return "E"  ;
    if (arc_index == 897) return "E"  ;
    if (arc_index == 898) return "E"  ;
    if (arc_index == 899) return "E"  ;
    if (arc_index == 900) return "E"  ;
    if (arc_index == 901) return "E"  ;
    if (arc_index == 907) return "E"  ;
    if (arc_index == 913) return "H"  ;
    if (arc_index == 950) return "H"  ;
    if (arc_index == 958) return "H"  ;
    if (arc_index == 963) return "H"  ;
    if (arc_index == 994) return "H"  ;
    if (arc_index == 1157) return "H"  ;
    if (arc_index == 1202) return "H"  ;
    if (arc_index == 1224) return "H"  ;
    if (arc_index == 1231) return "H"  ;
    if (arc_index == 1301) return "H"  ;
    if (arc_index == 1334) return "H"  ;
    if (arc_index == 1400) return "H"  ;
    if (arc_index == 1418) return "H"  ;
    if (arc_index == 1424) return "W"  ;
    if (arc_index == 1454) return "W"  ;
    if (arc_index == 1527) return "H"  ;
    if (arc_index == 1533) return "H"  ;
    if (arc_index == 1600) return "H"  ;
    if (arc_index == 1636) return "H"  ;
    if (arc_index == 1643) return "H"  ;
    if (arc_index == 1667) return "W"  ;
    if (arc_index == 1673) return "W"  ;
    if (arc_index == 1706) return "W"  ;
    if (arc_index == 1709) return "W"  ;
    if (arc_index == 1716) return "W"  ;
    if (arc_index == 1718) return "E"  ;
    if (arc_index == 1720) return "E"  ;
    if (arc_index == 1721) return "E"  ;
    if (arc_index == 1729) return "E"  ;
    if (arc_index == 1732) return "H"  ;
    if (arc_index == 1739) return "E"  ;
    if (arc_index == 1740) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1742) return "E"  ;
    if (arc_index == 1743) return "E"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1746) return "H"  ;
    if (arc_index == 1747) return "E"  ;
    if (arc_index == 1748) return "W"  ;
    if (arc_index == 1749) return "W"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1753) return "E"  ;
    if (arc_index == 1754) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1768) return "E"  ;
    if (arc_index == 1822) return "W"  ;
    if (arc_index == 1877) return "H"  ;
    if (arc_index == 1920) return "H"  ;
    if (arc_index == 1957) return "E"  ;
    if (arc_index == 1963) return "W"  ;
    if (arc_index == 1984) return "W"  ;
    if (arc_index == 1993) return "W"  ;
    if (arc_index == 2015) return "W"  ;
    if (arc_index == 2030) return "H"  ;
    if (arc_index == 2038) return "H"  ;
    if (arc_index == 2044) return "W"  ;
    if (arc_index == 2050) return "W"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2276) return "W"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2305) return "W"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2466) return "W"  ;
    if (arc_index == 2479) return "W"  ;
    if (arc_index == 2532) return "W"  ;
    if (arc_index == 2567) return "E"  ;
    if (arc_index == 2568) return "E"  ;
    if (arc_index == 2590) return "E"  ;
    if (arc_index == 2679) return "H"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2741) return "E"  ;
    if (arc_index == 2743) return "E"  ;
    if (arc_index == 2772) return "W"  ;
    if (arc_index == 2780) return "W"  ;
    if (arc_index == 2788) return "W"  ;
    if (arc_index == 2794) return "E"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2801) return "E"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2805) return "E"  ;
    if (arc_index == 2807) return "E"  ;
    if (arc_index == 2810) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2827) return "W"  ;
    if (arc_index == 2834) return "H"  ;
    if (arc_index == 2851) return "W"  ;
    if (arc_index == 2861) return "W"  ;
    if (arc_index == 2862) return "E"  ;
    if (arc_index == 2866) return "E"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2888) return "E"  ;
    if (arc_index == 2893) return "E"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 2)) begin 
    if (arc_index == 13) return "W"  ;
    if (arc_index == 63) return "H"  ;
    if (arc_index == 65) return "H"  ;
    if (arc_index == 71) return "H"  ;
    if (arc_index == 76) return "H"  ;
    if (arc_index == 79) return "H"  ;
    if (arc_index == 80) return "H"  ;
    if (arc_index == 106) return "H"  ;
    if (arc_index == 107) return "H"  ;
    if (arc_index == 115) return "H"  ;
    if (arc_index == 138) return "H"  ;
    if (arc_index == 148) return "W"  ;
    if (arc_index == 158) return "H"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 284) return "H"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 390) return "W"  ;
    if (arc_index == 395) return "H"  ;
    if (arc_index == 440) return "E"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 443) return "E"  ;
    if (arc_index == 454) return "E"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 456) return "E"  ;
    if (arc_index == 462) return "W"  ;
    if (arc_index == 465) return "H"  ;
    if (arc_index == 473) return "W"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 495) return "E"  ;
    if (arc_index == 501) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 520) return "E"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 591) return "E"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 640) return "H"  ;
    if (arc_index == 668) return "H"  ;
    if (arc_index == 687) return "H"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 751) return "W"  ;
    if (arc_index == 770) return "W"  ;
    if (arc_index == 779) return "W"  ;
    if (arc_index == 797) return "W"  ;
    if (arc_index == 799) return "W"  ;
    if (arc_index == 803) return "W"  ;
    if (arc_index == 808) return "W"  ;
    if (arc_index == 837) return "H"  ;
    if (arc_index == 865) return "H"  ;
    if (arc_index == 880) return "H"  ;
    if (arc_index == 886) return "W"  ;
    if (arc_index == 900) return "W"  ;
    if (arc_index == 902) return "W"  ;
    if (arc_index == 903) return "E"  ;
    if (arc_index == 904) return "E"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 906) return "E"  ;
    if (arc_index == 907) return "E"  ;
    if (arc_index == 908) return "E"  ;
    if (arc_index == 909) return "E"  ;
    if (arc_index == 910) return "E"  ;
    if (arc_index == 911) return "E"  ;
    if (arc_index == 912) return "E"  ;
    if (arc_index == 913) return "E"  ;
    if (arc_index == 914) return "E"  ;
    if (arc_index == 915) return "E"  ;
    if (arc_index == 916) return "E"  ;
    if (arc_index == 917) return "E"  ;
    if (arc_index == 918) return "E"  ;
    if (arc_index == 919) return "E"  ;
    if (arc_index == 920) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 923) return "E"  ;
    if (arc_index == 931) return "E"  ;
    if (arc_index == 935) return "H"  ;
    if (arc_index == 942) return "H"  ;
    if (arc_index == 946) return "H"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 980) return "H"  ;
    if (arc_index == 1010) return "H"  ;
    if (arc_index == 1017) return "E"  ;
    if (arc_index == 1063) return "E"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1179) return "H"  ;
    if (arc_index == 1190) return "E"  ;
    if (arc_index == 1191) return "E"  ;
    if (arc_index == 1192) return "E"  ;
    if (arc_index == 1193) return "E"  ;
    if (arc_index == 1197) return "E"  ;
    if (arc_index == 1202) return "E"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1208) return "E"  ;
    if (arc_index == 1209) return "E"  ;
    if (arc_index == 1213) return "E"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1225) return "E"  ;
    if (arc_index == 1231) return "E"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1356) return "H"  ;
    if (arc_index == 1366) return "H"  ;
    if (arc_index == 1438) return "H"  ;
    if (arc_index == 1440) return "H"  ;
    if (arc_index == 1465) return "H"  ;
    if (arc_index == 1466) return "H"  ;
    if (arc_index == 1503) return "H"  ;
    if (arc_index == 1527) return "H"  ;
    if (arc_index == 1533) return "H"  ;
    if (arc_index == 1549) return "H"  ;
    if (arc_index == 1563) return "H"  ;
    if (arc_index == 1605) return "E"  ;
    if (arc_index == 1634) return "W"  ;
    if (arc_index == 1637) return "W"  ;
    if (arc_index == 1642) return "W"  ;
    if (arc_index == 1644) return "W"  ;
    if (arc_index == 1664) return "W"  ;
    if (arc_index == 1665) return "H"  ;
    if (arc_index == 1690) return "W"  ;
    if (arc_index == 1715) return "W"  ;
    if (arc_index == 1719) return "W"  ;
    if (arc_index == 1723) return "W"  ;
    if (arc_index == 1726) return "W"  ;
    if (arc_index == 1735) return "W"  ;
    if (arc_index == 1740) return "W"  ;
    if (arc_index == 1743) return "W"  ;
    if (arc_index == 1752) return "W"  ;
    if (arc_index == 1754) return "H"  ;
    if (arc_index == 1768) return "H"  ;
    if (arc_index == 1785) return "W"  ;
    if (arc_index == 1790) return "W"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1823) return "W"  ;
    if (arc_index == 1831) return "W"  ;
    if (arc_index == 1835) return "W"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1899) return "H"  ;
    if (arc_index == 1921) return "H"  ;
    if (arc_index == 1929) return "H"  ;
    if (arc_index == 1931) return "E"  ;
    if (arc_index == 1935) return "E"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 1960) return "W"  ;
    if (arc_index == 2002) return "W"  ;
    if (arc_index == 2007) return "W"  ;
    if (arc_index == 2015) return "W"  ;
    if (arc_index == 2035) return "W"  ;
    if (arc_index == 2052) return "H"  ;
    if (arc_index == 2082) return "H"  ;
    if (arc_index == 2116) return "W"  ;
    if (arc_index == 2155) return "W"  ;
    if (arc_index == 2157) return "W"  ;
    if (arc_index == 2166) return "W"  ;
    if (arc_index == 2176) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2222) return "E"  ;
    if (arc_index == 2227) return "E"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2235) return "E"  ;
    if (arc_index == 2236) return "E"  ;
    if (arc_index == 2237) return "E"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2243) return "E"  ;
    if (arc_index == 2248) return "E"  ;
    if (arc_index == 2255) return "W"  ;
    if (arc_index == 2275) return "W"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2450) return "W"  ;
    if (arc_index == 2452) return "W"  ;
    if (arc_index == 2469) return "W"  ;
    if (arc_index == 2485) return "W"  ;
    if (arc_index == 2526) return "W"  ;
    if (arc_index == 2555) return "W"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2576) return "E"  ;
    if (arc_index == 2589) return "E"  ;
    if (arc_index == 2590) return "E"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2662) return "E"  ;
    if (arc_index == 2664) return "E"  ;
    if (arc_index == 2669) return "E"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2677) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2701) return "H"  ;
    if (arc_index == 2730) return "H"  ;
    if (arc_index == 2733) return "H"  ;
    if (arc_index == 2746) return "H"  ;
    if (arc_index == 2765) return "H"  ;
    if (arc_index == 2796) return "E"  ;
    if (arc_index == 2812) return "E"  ;
    if (arc_index == 2856) return "H"  ;
    if (arc_index == 2868) return "H"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 2)) begin 
    if (arc_index == 67) return "E"  ;
    if (arc_index == 73) return "E"  ;
    if (arc_index == 85) return "H"  ;
    if (arc_index == 93) return "H"  ;
    if (arc_index == 99) return "H"  ;
    if (arc_index == 112) return "W"  ;
    if (arc_index == 115) return "W"  ;
    if (arc_index == 135) return "W"  ;
    if (arc_index == 144) return "W"  ;
    if (arc_index == 145) return "W"  ;
    if (arc_index == 180) return "H"  ;
    if (arc_index == 285) return "H"  ;
    if (arc_index == 306) return "H"  ;
    if (arc_index == 352) return "W"  ;
    if (arc_index == 357) return "W"  ;
    if (arc_index == 374) return "E"  ;
    if (arc_index == 376) return "E"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 382) return "E"  ;
    if (arc_index == 385) return "E"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 387) return "E"  ;
    if (arc_index == 392) return "E"  ;
    if (arc_index == 393) return "E"  ;
    if (arc_index == 417) return "H"  ;
    if (arc_index == 451) return "E"  ;
    if (arc_index == 487) return "H"  ;
    if (arc_index == 513) return "H"  ;
    if (arc_index == 530) return "H"  ;
    if (arc_index == 641) return "H"  ;
    if (arc_index == 651) return "W"  ;
    if (arc_index == 662) return "H"  ;
    if (arc_index == 679) return "H"  ;
    if (arc_index == 681) return "H"  ;
    if (arc_index == 770) return "H"  ;
    if (arc_index == 792) return "H"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 797) return "E"  ;
    if (arc_index == 799) return "E"  ;
    if (arc_index == 800) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 803) return "E"  ;
    if (arc_index == 807) return "E"  ;
    if (arc_index == 808) return "E"  ;
    if (arc_index == 809) return "E"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 811) return "E"  ;
    if (arc_index == 812) return "E"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 859) return "H"  ;
    if (arc_index == 865) return "H"  ;
    if (arc_index == 902) return "H"  ;
    if (arc_index == 924) return "H"  ;
    if (arc_index == 925) return "H"  ;
    if (arc_index == 926) return "H"  ;
    if (arc_index == 927) return "H"  ;
    if (arc_index == 928) return "H"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 931) return "E"  ;
    if (arc_index == 932) return "E"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 934) return "E"  ;
    if (arc_index == 935) return "E"  ;
    if (arc_index == 936) return "E"  ;
    if (arc_index == 937) return "E"  ;
    if (arc_index == 938) return "E"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 940) return "E"  ;
    if (arc_index == 941) return "E"  ;
    if (arc_index == 942) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 957) return "H"  ;
    if (arc_index == 1002) return "H"  ;
    if (arc_index == 1011) return "H"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1032) return "E"  ;
    if (arc_index == 1123) return "E"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1201) return "H"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1240) return "W"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1371) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1378) return "H"  ;
    if (arc_index == 1462) return "H"  ;
    if (arc_index == 1496) return "H"  ;
    if (arc_index == 1528) return "H"  ;
    if (arc_index == 1529) return "E"  ;
    if (arc_index == 1536) return "E"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1571) return "H"  ;
    if (arc_index == 1603) return "E"  ;
    if (arc_index == 1644) return "E"  ;
    if (arc_index == 1658) return "E"  ;
    if (arc_index == 1687) return "H"  ;
    if (arc_index == 1740) return "H"  ;
    if (arc_index == 1743) return "W"  ;
    if (arc_index == 1776) return "H"  ;
    if (arc_index == 1789) return "H"  ;
    if (arc_index == 1790) return "H"  ;
    if (arc_index == 1864) return "W"  ;
    if (arc_index == 1878) return "W"  ;
    if (arc_index == 1921) return "H"  ;
    if (arc_index == 1935) return "E"  ;
    if (arc_index == 1937) return "E"  ;
    if (arc_index == 1942) return "E"  ;
    if (arc_index == 2002) return "E"  ;
    if (arc_index == 2004) return "E"  ;
    if (arc_index == 2006) return "E"  ;
    if (arc_index == 2007) return "E"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2013) return "E"  ;
    if (arc_index == 2014) return "E"  ;
    if (arc_index == 2015) return "E"  ;
    if (arc_index == 2020) return "E"  ;
    if (arc_index == 2021) return "E"  ;
    if (arc_index == 2023) return "E"  ;
    if (arc_index == 2035) return "E"  ;
    if (arc_index == 2074) return "H"  ;
    if (arc_index == 2162) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2461) return "W"  ;
    if (arc_index == 2515) return "W"  ;
    if (arc_index == 2526) return "W"  ;
    if (arc_index == 2527) return "W"  ;
    if (arc_index == 2584) return "W"  ;
    if (arc_index == 2586) return "E"  ;
    if (arc_index == 2588) return "E"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2723) return "H"  ;
    if (arc_index == 2746) return "H"  ;
    if (arc_index == 2747) return "H"  ;
    if (arc_index == 2765) return "H"  ;
    if (arc_index == 2854) return "H"  ;
    if (arc_index == 2868) return "H"  ;
    if (arc_index == 2878) return "H"  ;
    if (arc_index == 2879) return "H"  ;
    if (arc_index == 2887) return "H"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 0)) begin 
    if (arc_index == 107) return "H"  ;
    if (arc_index == 115) return "H"  ;
    if (arc_index == 202) return "H"  ;
    if (arc_index == 328) return "H"  ;
    if (arc_index == 388) return "H"  ;
    if (arc_index == 439) return "H"  ;
    if (arc_index == 492) return "H"  ;
    if (arc_index == 493) return "E"  ;
    if (arc_index == 509) return "H"  ;
    if (arc_index == 577) return "E"  ;
    if (arc_index == 581) return "E"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 587) return "E"  ;
    if (arc_index == 684) return "H"  ;
    if (arc_index == 761) return "H"  ;
    if (arc_index == 800) return "H"  ;
    if (arc_index == 849) return "H"  ;
    if (arc_index == 881) return "H"  ;
    if (arc_index == 924) return "H"  ;
    if (arc_index == 931) return "H"  ;
    if (arc_index == 946) return "E"  ;
    if (arc_index == 947) return "E"  ;
    if (arc_index == 948) return "E"  ;
    if (arc_index == 949) return "E"  ;
    if (arc_index == 950) return "E"  ;
    if (arc_index == 951) return "E"  ;
    if (arc_index == 952) return "E"  ;
    if (arc_index == 953) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 957) return "E"  ;
    if (arc_index == 958) return "E"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 960) return "E"  ;
    if (arc_index == 961) return "E"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 964) return "E"  ;
    if (arc_index == 965) return "E"  ;
    if (arc_index == 966) return "E"  ;
    if (arc_index == 967) return "E"  ;
    if (arc_index == 979) return "H"  ;
    if (arc_index == 1024) return "H"  ;
    if (arc_index == 1223) return "H"  ;
    if (arc_index == 1400) return "H"  ;
    if (arc_index == 1424) return "H"  ;
    if (arc_index == 1484) return "H"  ;
    if (arc_index == 1593) return "H"  ;
    if (arc_index == 1601) return "E"  ;
    if (arc_index == 1709) return "H"  ;
    if (arc_index == 1722) return "H"  ;
    if (arc_index == 1733) return "H"  ;
    if (arc_index == 1798) return "H"  ;
    if (arc_index == 1812) return "H"  ;
    if (arc_index == 1943) return "H"  ;
    if (arc_index == 2021) return "H"  ;
    if (arc_index == 2044) return "H"  ;
    if (arc_index == 2096) return "H"  ;
    if (arc_index == 2116) return "H"  ;
    if (arc_index == 2242) return "H"  ;
    if (arc_index == 2423) return "H"  ;
    if (arc_index == 2663) return "H"  ;
    if (arc_index == 2671) return "H"  ;
    if (arc_index == 2734) return "H"  ;
    if (arc_index == 2740) return "H"  ;
    if (arc_index == 2745) return "H"  ;
    if (arc_index == 2860) return "H"  ;
    if (arc_index == 2863) return "H"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2868) return "E"  ;
    if (arc_index == 2869) return "E"  ;
    if (arc_index == 2874) return "E"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2879) return "E"  ;
    if (arc_index == 2880) return "E"  ;
    if (arc_index == 2881) return "E"  ;
    if (arc_index == 2900) return "H"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 5)) begin 
    if (arc_index == 0) return "W"  ;
    if (arc_index == 23) return "W"  ;
    if (arc_index == 24) return "E"  ;
    if (arc_index == 29) return "E"  ;
    if (arc_index == 30) return "E"  ;
    if (arc_index == 31) return "E"  ;
    if (arc_index == 33) return "E"  ;
    if (arc_index == 37) return "E"  ;
    if (arc_index == 39) return "E"  ;
    if (arc_index == 43) return "E"  ;
    if (arc_index == 100) return "W"  ;
    if (arc_index == 106) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 113) return "E"  ;
    if (arc_index == 116) return "E"  ;
    if (arc_index == 117) return "W"  ;
    if (arc_index == 118) return "E"  ;
    if (arc_index == 119) return "E"  ;
    if (arc_index == 122) return "W"  ;
    if (arc_index == 123) return "W"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 125) return "E"  ;
    if (arc_index == 128) return "E"  ;
    if (arc_index == 129) return "H"  ;
    if (arc_index == 130) return "H"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 137) return "H"  ;
    if (arc_index == 149) return "E"  ;
    if (arc_index == 163) return "E"  ;
    if (arc_index == 165) return "E"  ;
    if (arc_index == 180) return "W"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 210) return "W"  ;
    if (arc_index == 224) return "H"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 229) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 279) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 299) return "W"  ;
    if (arc_index == 345) return "W"  ;
    if (arc_index == 350) return "H"  ;
    if (arc_index == 362) return "H"  ;
    if (arc_index == 366) return "H"  ;
    if (arc_index == 367) return "H"  ;
    if (arc_index == 371) return "W"  ;
    if (arc_index == 377) return "W"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 399) return "E"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 404) return "W"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 412) return "W"  ;
    if (arc_index == 414) return "W"  ;
    if (arc_index == 445) return "E"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 461) return "H"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 474) return "E"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 531) return "H"  ;
    if (arc_index == 640) return "W"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 706) return "H"  ;
    if (arc_index == 726) return "H"  ;
    if (arc_index == 734) return "H"  ;
    if (arc_index == 739) return "H"  ;
    if (arc_index == 757) return "H"  ;
    if (arc_index == 759) return "E"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 828) return "E"  ;
    if (arc_index == 850) return "E"  ;
    if (arc_index == 862) return "E"  ;
    if (arc_index == 874) return "W"  ;
    if (arc_index == 879) return "W"  ;
    if (arc_index == 891) return "W"  ;
    if (arc_index == 903) return "H"  ;
    if (arc_index == 929) return "H"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 946) return "H"  ;
    if (arc_index == 962) return "H"  ;
    if (arc_index == 968) return "H"  ;
    if (arc_index == 969) return "E"  ;
    if (arc_index == 970) return "E"  ;
    if (arc_index == 971) return "E"  ;
    if (arc_index == 972) return "E"  ;
    if (arc_index == 973) return "E"  ;
    if (arc_index == 974) return "E"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 976) return "E"  ;
    if (arc_index == 977) return "E"  ;
    if (arc_index == 978) return "W"  ;
    if (arc_index == 979) return "W"  ;
    if (arc_index == 980) return "W"  ;
    if (arc_index == 981) return "W"  ;
    if (arc_index == 982) return "E"  ;
    if (arc_index == 983) return "E"  ;
    if (arc_index == 984) return "E"  ;
    if (arc_index == 985) return "E"  ;
    if (arc_index == 986) return "E"  ;
    if (arc_index == 987) return "E"  ;
    if (arc_index == 988) return "E"  ;
    if (arc_index == 989) return "E"  ;
    if (arc_index == 991) return "E"  ;
    if (arc_index == 993) return "E"  ;
    if (arc_index == 997) return "E"  ;
    if (arc_index == 1001) return "H"  ;
    if (arc_index == 1006) return "H"  ;
    if (arc_index == 1014) return "E"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1046) return "H"  ;
    if (arc_index == 1059) return "H"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1166) return "W"  ;
    if (arc_index == 1169) return "W"  ;
    if (arc_index == 1172) return "W"  ;
    if (arc_index == 1179) return "W"  ;
    if (arc_index == 1184) return "W"  ;
    if (arc_index == 1189) return "E"  ;
    if (arc_index == 1199) return "E"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1211) return "E"  ;
    if (arc_index == 1217) return "E"  ;
    if (arc_index == 1218) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1245) return "H"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1266) return "W"  ;
    if (arc_index == 1288) return "W"  ;
    if (arc_index == 1289) return "W"  ;
    if (arc_index == 1293) return "W"  ;
    if (arc_index == 1295) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1365) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1393) return "W"  ;
    if (arc_index == 1422) return "H"  ;
    if (arc_index == 1431) return "H"  ;
    if (arc_index == 1433) return "E"  ;
    if (arc_index == 1439) return "W"  ;
    if (arc_index == 1442) return "E"  ;
    if (arc_index == 1447) return "E"  ;
    if (arc_index == 1470) return "W"  ;
    if (arc_index == 1498) return "W"  ;
    if (arc_index == 1499) return "W"  ;
    if (arc_index == 1500) return "E"  ;
    if (arc_index == 1506) return "H"  ;
    if (arc_index == 1507) return "E"  ;
    if (arc_index == 1508) return "E"  ;
    if (arc_index == 1514) return "E"  ;
    if (arc_index == 1515) return "E"  ;
    if (arc_index == 1517) return "E"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1522) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1546) return "E"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1592) return "W"  ;
    if (arc_index == 1615) return "H"  ;
    if (arc_index == 1621) return "H"  ;
    if (arc_index == 1635) return "H"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1710) return "E"  ;
    if (arc_index == 1731) return "H"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1773) return "E"  ;
    if (arc_index == 1820) return "H"  ;
    if (arc_index == 1821) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1834) return "H"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1855) return "E"  ;
    if (arc_index == 1872) return "E"  ;
    if (arc_index == 1881) return "E"  ;
    if (arc_index == 1883) return "E"  ;
    if (arc_index == 1884) return "E"  ;
    if (arc_index == 1902) return "E"  ;
    if (arc_index == 1909) return "E"  ;
    if (arc_index == 1923) return "E"  ;
    if (arc_index == 1929) return "E"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 1965) return "H"  ;
    if (arc_index == 1973) return "W"  ;
    if (arc_index == 1976) return "W"  ;
    if (arc_index == 2004) return "W"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2061) return "E"  ;
    if (arc_index == 2064) return "E"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2112) return "W"  ;
    if (arc_index == 2117) return "W"  ;
    if (arc_index == 2118) return "H"  ;
    if (arc_index == 2119) return "H"  ;
    if (arc_index == 2130) return "E"  ;
    if (arc_index == 2141) return "E"  ;
    if (arc_index == 2163) return "E"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2202) return "W"  ;
    if (arc_index == 2204) return "W"  ;
    if (arc_index == 2229) return "W"  ;
    if (arc_index == 2259) return "W"  ;
    if (arc_index == 2279) return "W"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2330) return "W"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2398) return "W"  ;
    if (arc_index == 2426) return "E"  ;
    if (arc_index == 2427) return "E"  ;
    if (arc_index == 2428) return "E"  ;
    if (arc_index == 2430) return "E"  ;
    if (arc_index == 2431) return "E"  ;
    if (arc_index == 2435) return "E"  ;
    if (arc_index == 2439) return "E"  ;
    if (arc_index == 2449) return "E"  ;
    if (arc_index == 2491) return "E"  ;
    if (arc_index == 2493) return "E"  ;
    if (arc_index == 2498) return "W"  ;
    if (arc_index == 2521) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2524) return "E"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2704) return "E"  ;
    if (arc_index == 2767) return "H"  ;
    if (arc_index == 2771) return "E"  ;
    if (arc_index == 2774) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2922) return "H"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 3)) begin 
    if (arc_index == 18) return "H"  ;
    if (arc_index == 42) return "H"  ;
    if (arc_index == 48) return "W"  ;
    if (arc_index == 102) return "W"  ;
    if (arc_index == 141) return "W"  ;
    if (arc_index == 144) return "W"  ;
    if (arc_index == 151) return "H"  ;
    if (arc_index == 159) return "H"  ;
    if (arc_index == 173) return "H"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 246) return "H"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 355) return "W"  ;
    if (arc_index == 372) return "H"  ;
    if (arc_index == 392) return "E"  ;
    if (arc_index == 418) return "W"  ;
    if (arc_index == 434) return "W"  ;
    if (arc_index == 483) return "H"  ;
    if (arc_index == 513) return "E"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 553) return "H"  ;
    if (arc_index == 586) return "H"  ;
    if (arc_index == 638) return "H"  ;
    if (arc_index == 645) return "W"  ;
    if (arc_index == 663) return "W"  ;
    if (arc_index == 664) return "W"  ;
    if (arc_index == 666) return "E"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 668) return "E"  ;
    if (arc_index == 674) return "E"  ;
    if (arc_index == 675) return "E"  ;
    if (arc_index == 676) return "E"  ;
    if (arc_index == 678) return "E"  ;
    if (arc_index == 679) return "E"  ;
    if (arc_index == 693) return "E"  ;
    if (arc_index == 727) return "W"  ;
    if (arc_index == 728) return "H"  ;
    if (arc_index == 732) return "H"  ;
    if (arc_index == 793) return "E"  ;
    if (arc_index == 795) return "E"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 804) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 806) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 825) return "W"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 870) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 925) return "H"  ;
    if (arc_index == 927) return "E"  ;
    if (arc_index == 937) return "E"  ;
    if (arc_index == 968) return "H"  ;
    if (arc_index == 990) return "H"  ;
    if (arc_index == 991) return "E"  ;
    if (arc_index == 992) return "E"  ;
    if (arc_index == 993) return "E"  ;
    if (arc_index == 994) return "E"  ;
    if (arc_index == 995) return "E"  ;
    if (arc_index == 996) return "E"  ;
    if (arc_index == 997) return "E"  ;
    if (arc_index == 998) return "E"  ;
    if (arc_index == 999) return "E"  ;
    if (arc_index == 1000) return "E"  ;
    if (arc_index == 1001) return "E"  ;
    if (arc_index == 1002) return "E"  ;
    if (arc_index == 1003) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1007) return "E"  ;
    if (arc_index == 1008) return "E"  ;
    if (arc_index == 1009) return "E"  ;
    if (arc_index == 1010) return "E"  ;
    if (arc_index == 1011) return "W"  ;
    if (arc_index == 1014) return "W"  ;
    if (arc_index == 1019) return "E"  ;
    if (arc_index == 1023) return "H"  ;
    if (arc_index == 1033) return "H"  ;
    if (arc_index == 1068) return "H"  ;
    if (arc_index == 1069) return "W"  ;
    if (arc_index == 1123) return "W"  ;
    if (arc_index == 1198) return "W"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1246) return "W"  ;
    if (arc_index == 1267) return "H"  ;
    if (arc_index == 1289) return "H"  ;
    if (arc_index == 1371) return "H"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1381) return "W"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1439) return "W"  ;
    if (arc_index == 1444) return "H"  ;
    if (arc_index == 1447) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1496) return "W"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1528) return "H"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1637) return "H"  ;
    if (arc_index == 1657) return "H"  ;
    if (arc_index == 1753) return "H"  ;
    if (arc_index == 1775) return "H"  ;
    if (arc_index == 1842) return "H"  ;
    if (arc_index == 1856) return "H"  ;
    if (arc_index == 1987) return "H"  ;
    if (arc_index == 2017) return "E"  ;
    if (arc_index == 2067) return "W"  ;
    if (arc_index == 2137) return "W"  ;
    if (arc_index == 2140) return "H"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2440) return "W"  ;
    if (arc_index == 2442) return "W"  ;
    if (arc_index == 2443) return "W"  ;
    if (arc_index == 2450) return "W"  ;
    if (arc_index == 2453) return "W"  ;
    if (arc_index == 2456) return "W"  ;
    if (arc_index == 2461) return "W"  ;
    if (arc_index == 2509) return "W"  ;
    if (arc_index == 2513) return "E"  ;
    if (arc_index == 2514) return "E"  ;
    if (arc_index == 2520) return "E"  ;
    if (arc_index == 2540) return "E"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2577) return "E"  ;
    if (arc_index == 2578) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2592) return "E"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2747) return "W"  ;
    if (arc_index == 2755) return "W"  ;
    if (arc_index == 2789) return "H"  ;
    if (arc_index == 2842) return "H"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 1)) begin 
    if (arc_index == 40) return "H"  ;
    if (arc_index == 173) return "H"  ;
    if (arc_index == 181) return "H"  ;
    if (arc_index == 268) return "H"  ;
    if (arc_index == 394) return "H"  ;
    if (arc_index == 407) return "H"  ;
    if (arc_index == 505) return "H"  ;
    if (arc_index == 575) return "H"  ;
    if (arc_index == 750) return "H"  ;
    if (arc_index == 947) return "H"  ;
    if (arc_index == 990) return "H"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1013) return "E"  ;
    if (arc_index == 1014) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1017) return "E"  ;
    if (arc_index == 1018) return "E"  ;
    if (arc_index == 1019) return "E"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1021) return "E"  ;
    if (arc_index == 1022) return "E"  ;
    if (arc_index == 1023) return "E"  ;
    if (arc_index == 1024) return "E"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1026) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1029) return "E"  ;
    if (arc_index == 1030) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1032) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1045) return "H"  ;
    if (arc_index == 1090) return "H"  ;
    if (arc_index == 1289) return "H"  ;
    if (arc_index == 1466) return "H"  ;
    if (arc_index == 1526) return "E"  ;
    if (arc_index == 1550) return "H"  ;
    if (arc_index == 1659) return "H"  ;
    if (arc_index == 1775) return "H"  ;
    if (arc_index == 1864) return "H"  ;
    if (arc_index == 1878) return "H"  ;
    if (arc_index == 2009) return "H"  ;
    if (arc_index == 2162) return "H"  ;
    if (arc_index == 2811) return "H"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 11)) begin 
    if (arc_index == 62) return "H"  ;
    if (arc_index == 168) return "H"  ;
    if (arc_index == 195) return "H"  ;
    if (arc_index == 203) return "H"  ;
    if (arc_index == 290) return "H"  ;
    if (arc_index == 416) return "H"  ;
    if (arc_index == 477) return "H"  ;
    if (arc_index == 527) return "H"  ;
    if (arc_index == 566) return "H"  ;
    if (arc_index == 580) return "H"  ;
    if (arc_index == 597) return "H"  ;
    if (arc_index == 711) return "H"  ;
    if (arc_index == 772) return "H"  ;
    if (arc_index == 969) return "H"  ;
    if (arc_index == 1012) return "H"  ;
    if (arc_index == 1034) return "H"  ;
    if (arc_index == 1035) return "W"  ;
    if (arc_index == 1036) return "W"  ;
    if (arc_index == 1037) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1039) return "W"  ;
    if (arc_index == 1040) return "W"  ;
    if (arc_index == 1041) return "W"  ;
    if (arc_index == 1042) return "W"  ;
    if (arc_index == 1043) return "W"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1046) return "W"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1048) return "W"  ;
    if (arc_index == 1049) return "W"  ;
    if (arc_index == 1050) return "W"  ;
    if (arc_index == 1051) return "W"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1053) return "W"  ;
    if (arc_index == 1054) return "W"  ;
    if (arc_index == 1055) return "W"  ;
    if (arc_index == 1067) return "H"  ;
    if (arc_index == 1112) return "H"  ;
    if (arc_index == 1311) return "H"  ;
    if (arc_index == 1488) return "H"  ;
    if (arc_index == 1572) return "H"  ;
    if (arc_index == 1573) return "H"  ;
    if (arc_index == 1668) return "H"  ;
    if (arc_index == 1681) return "H"  ;
    if (arc_index == 1797) return "H"  ;
    if (arc_index == 1809) return "H"  ;
    if (arc_index == 1886) return "H"  ;
    if (arc_index == 1900) return "H"  ;
    if (arc_index == 2031) return "H"  ;
    if (arc_index == 2133) return "H"  ;
    if (arc_index == 2184) return "H"  ;
    if (arc_index == 2203) return "H"  ;
    if (arc_index == 2378) return "H"  ;
    if (arc_index == 2618) return "H"  ;
    if (arc_index == 2641) return "H"  ;
    if (arc_index == 2642) return "H"  ;
    if (arc_index == 2643) return "H"  ;
    if (arc_index == 2644) return "H"  ;
    if (arc_index == 2645) return "H"  ;
    if (arc_index == 2647) return "H"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2651) return "W"  ;
    if (arc_index == 2653) return "W"  ;
    if (arc_index == 2654) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2658) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2718) return "W"  ;
    if (arc_index == 2726) return "W"  ;
    if (arc_index == 2833) return "H"  ;
    if (arc_index == 2917) return "H"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 7)) begin 
    if (arc_index == 2) return "E"  ;
    if (arc_index == 8) return "E"  ;
    if (arc_index == 10) return "E"  ;
    if (arc_index == 11) return "E"  ;
    if (arc_index == 15) return "E"  ;
    if (arc_index == 17) return "E"  ;
    if (arc_index == 21) return "E"  ;
    if (arc_index == 43) return "E"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 84) return "H"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 92) return "E"  ;
    if (arc_index == 95) return "E"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 156) return "E"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 165) return "W"  ;
    if (arc_index == 170) return "W"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 176) return "W"  ;
    if (arc_index == 198) return "E"  ;
    if (arc_index == 201) return "E"  ;
    if (arc_index == 206) return "E"  ;
    if (arc_index == 209) return "E"  ;
    if (arc_index == 217) return "H"  ;
    if (arc_index == 219) return "E"  ;
    if (arc_index == 225) return "H"  ;
    if (arc_index == 233) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 265) return "W"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 269) return "W"  ;
    if (arc_index == 270) return "W"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 277) return "W"  ;
    if (arc_index == 284) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 296) return "W"  ;
    if (arc_index == 308) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 312) return "H"  ;
    if (arc_index == 315) return "W"  ;
    if (arc_index == 332) return "E"  ;
    if (arc_index == 342) return "E"  ;
    if (arc_index == 344) return "E"  ;
    if (arc_index == 347) return "E"  ;
    if (arc_index == 354) return "E"  ;
    if (arc_index == 359) return "E"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 428) return "E"  ;
    if (arc_index == 433) return "E"  ;
    if (arc_index == 438) return "H"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 481) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 537) return "E"  ;
    if (arc_index == 538) return "W"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 549) return "H"  ;
    if (arc_index == 554) return "H"  ;
    if (arc_index == 561) return "H"  ;
    if (arc_index == 564) return "H"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 595) return "E"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 603) return "W"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 607) return "W"  ;
    if (arc_index == 609) return "W"  ;
    if (arc_index == 610) return "W"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 619) return "H"  ;
    if (arc_index == 643) return "E"  ;
    if (arc_index == 652) return "E"  ;
    if (arc_index == 653) return "E"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 677) return "E"  ;
    if (arc_index == 695) return "E"  ;
    if (arc_index == 703) return "E"  ;
    if (arc_index == 713) return "E"  ;
    if (arc_index == 736) return "E"  ;
    if (arc_index == 742) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 794) return "H"  ;
    if (arc_index == 828) return "H"  ;
    if (arc_index == 829) return "H"  ;
    if (arc_index == 831) return "H"  ;
    if (arc_index == 857) return "H"  ;
    if (arc_index == 917) return "E"  ;
    if (arc_index == 973) return "E"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 991) return "H"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1034) return "H"  ;
    if (arc_index == 1035) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1056) return "W"  ;
    if (arc_index == 1057) return "W"  ;
    if (arc_index == 1058) return "E"  ;
    if (arc_index == 1059) return "E"  ;
    if (arc_index == 1060) return "E"  ;
    if (arc_index == 1061) return "W"  ;
    if (arc_index == 1062) return "W"  ;
    if (arc_index == 1063) return "W"  ;
    if (arc_index == 1064) return "W"  ;
    if (arc_index == 1065) return "W"  ;
    if (arc_index == 1066) return "E"  ;
    if (arc_index == 1067) return "E"  ;
    if (arc_index == 1068) return "W"  ;
    if (arc_index == 1069) return "W"  ;
    if (arc_index == 1070) return "W"  ;
    if (arc_index == 1071) return "E"  ;
    if (arc_index == 1072) return "E"  ;
    if (arc_index == 1073) return "E"  ;
    if (arc_index == 1074) return "E"  ;
    if (arc_index == 1075) return "W"  ;
    if (arc_index == 1076) return "W"  ;
    if (arc_index == 1077) return "W"  ;
    if (arc_index == 1086) return "W"  ;
    if (arc_index == 1089) return "H"  ;
    if (arc_index == 1116) return "E"  ;
    if (arc_index == 1119) return "E"  ;
    if (arc_index == 1133) return "W"  ;
    if (arc_index == 1134) return "H"  ;
    if (arc_index == 1144) return "H"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1148) return "W"  ;
    if (arc_index == 1150) return "W"  ;
    if (arc_index == 1177) return "E"  ;
    if (arc_index == 1186) return "E"  ;
    if (arc_index == 1274) return "W"  ;
    if (arc_index == 1280) return "W"  ;
    if (arc_index == 1286) return "W"  ;
    if (arc_index == 1290) return "W"  ;
    if (arc_index == 1297) return "W"  ;
    if (arc_index == 1313) return "W"  ;
    if (arc_index == 1321) return "W"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1325) return "W"  ;
    if (arc_index == 1327) return "W"  ;
    if (arc_index == 1328) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1333) return "H"  ;
    if (arc_index == 1334) return "H"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1367) return "W"  ;
    if (arc_index == 1374) return "W"  ;
    if (arc_index == 1375) return "E"  ;
    if (arc_index == 1379) return "E"  ;
    if (arc_index == 1427) return "E"  ;
    if (arc_index == 1445) return "E"  ;
    if (arc_index == 1480) return "W"  ;
    if (arc_index == 1490) return "W"  ;
    if (arc_index == 1494) return "W"  ;
    if (arc_index == 1507) return "E"  ;
    if (arc_index == 1510) return "H"  ;
    if (arc_index == 1515) return "H"  ;
    if (arc_index == 1541) return "H"  ;
    if (arc_index == 1542) return "H"  ;
    if (arc_index == 1543) return "H"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1594) return "H"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1672) return "W"  ;
    if (arc_index == 1673) return "W"  ;
    if (arc_index == 1689) return "W"  ;
    if (arc_index == 1696) return "W"  ;
    if (arc_index == 1703) return "H"  ;
    if (arc_index == 1734) return "H"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1764) return "E"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1803) return "E"  ;
    if (arc_index == 1807) return "W"  ;
    if (arc_index == 1810) return "W"  ;
    if (arc_index == 1813) return "W"  ;
    if (arc_index == 1814) return "W"  ;
    if (arc_index == 1818) return "W"  ;
    if (arc_index == 1819) return "H"  ;
    if (arc_index == 1820) return "H"  ;
    if (arc_index == 1821) return "H"  ;
    if (arc_index == 1823) return "W"  ;
    if (arc_index == 1829) return "W"  ;
    if (arc_index == 1836) return "W"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1893) return "W"  ;
    if (arc_index == 1901) return "W"  ;
    if (arc_index == 1903) return "E"  ;
    if (arc_index == 1907) return "E"  ;
    if (arc_index == 1908) return "H"  ;
    if (arc_index == 1922) return "H"  ;
    if (arc_index == 1936) return "H"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1953) return "E"  ;
    if (arc_index == 1958) return "E"  ;
    if (arc_index == 1959) return "E"  ;
    if (arc_index == 1963) return "E"  ;
    if (arc_index == 1966) return "W"  ;
    if (arc_index == 1971) return "W"  ;
    if (arc_index == 1977) return "W"  ;
    if (arc_index == 1978) return "W"  ;
    if (arc_index == 1979) return "W"  ;
    if (arc_index == 1991) return "W"  ;
    if (arc_index == 1994) return "W"  ;
    if (arc_index == 2036) return "W"  ;
    if (arc_index == 2042) return "W"  ;
    if (arc_index == 2053) return "H"  ;
    if (arc_index == 2075) return "H"  ;
    if (arc_index == 2087) return "W"  ;
    if (arc_index == 2159) return "W"  ;
    if (arc_index == 2182) return "W"  ;
    if (arc_index == 2206) return "H"  ;
    if (arc_index == 2215) return "H"  ;
    if (arc_index == 2249) return "E"  ;
    if (arc_index == 2258) return "E"  ;
    if (arc_index == 2266) return "E"  ;
    if (arc_index == 2268) return "E"  ;
    if (arc_index == 2285) return "E"  ;
    if (arc_index == 2286) return "E"  ;
    if (arc_index == 2287) return "E"  ;
    if (arc_index == 2288) return "E"  ;
    if (arc_index == 2296) return "E"  ;
    if (arc_index == 2299) return "E"  ;
    if (arc_index == 2306) return "E"  ;
    if (arc_index == 2318) return "E"  ;
    if (arc_index == 2320) return "W"  ;
    if (arc_index == 2321) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2386) return "W"  ;
    if (arc_index == 2389) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2413) return "W"  ;
    if (arc_index == 2419) return "W"  ;
    if (arc_index == 2432) return "W"  ;
    if (arc_index == 2451) return "W"  ;
    if (arc_index == 2496) return "W"  ;
    if (arc_index == 2507) return "W"  ;
    if (arc_index == 2523) return "W"  ;
    if (arc_index == 2537) return "E"  ;
    if (arc_index == 2538) return "E"  ;
    if (arc_index == 2543) return "E"  ;
    if (arc_index == 2548) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2605) return "E"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2620) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2670) return "W"  ;
    if (arc_index == 2684) return "W"  ;
    if (arc_index == 2689) return "E"  ;
    if (arc_index == 2690) return "E"  ;
    if (arc_index == 2696) return "E"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2714) return "W"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2810) return "E"  ;
    if (arc_index == 2819) return "E"  ;
    if (arc_index == 2820) return "E"  ;
    if (arc_index == 2821) return "E"  ;
    if (arc_index == 2824) return "E"  ;
    if (arc_index == 2825) return "E"  ;
    if (arc_index == 2837) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2855) return "H"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2895) return "E"  ;
    if (arc_index == 2902) return "E"  ;
    if (arc_index == 2904) return "W"  ;
    if (arc_index == 2912) return "W"  ;
    if (arc_index == 2915) return "W"  ;
    if (arc_index == 2922) return "W"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 1)) begin 
    if (arc_index == 79) return "W"  ;
    if (arc_index == 106) return "H"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 115) return "W"  ;
    if (arc_index == 145) return "W"  ;
    if (arc_index == 202) return "W"  ;
    if (arc_index == 239) return "H"  ;
    if (arc_index == 244) return "H"  ;
    if (arc_index == 247) return "H"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 334) return "H"  ;
    if (arc_index == 389) return "H"  ;
    if (arc_index == 406) return "H"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 449) return "W"  ;
    if (arc_index == 450) return "W"  ;
    if (arc_index == 460) return "H"  ;
    if (arc_index == 478) return "H"  ;
    if (arc_index == 486) return "H"  ;
    if (arc_index == 493) return "H"  ;
    if (arc_index == 508) return "H"  ;
    if (arc_index == 515) return "H"  ;
    if (arc_index == 550) return "H"  ;
    if (arc_index == 571) return "H"  ;
    if (arc_index == 577) return "E"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 587) return "E"  ;
    if (arc_index == 641) return "H"  ;
    if (arc_index == 654) return "H"  ;
    if (arc_index == 668) return "H"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 753) return "W"  ;
    if (arc_index == 761) return "W"  ;
    if (arc_index == 773) return "W"  ;
    if (arc_index == 774) return "W"  ;
    if (arc_index == 783) return "W"  ;
    if (arc_index == 799) return "W"  ;
    if (arc_index == 800) return "W"  ;
    if (arc_index == 816) return "H"  ;
    if (arc_index == 894) return "H"  ;
    if (arc_index == 931) return "W"  ;
    if (arc_index == 946) return "W"  ;
    if (arc_index == 948) return "W"  ;
    if (arc_index == 949) return "E"  ;
    if (arc_index == 950) return "E"  ;
    if (arc_index == 951) return "E"  ;
    if (arc_index == 952) return "E"  ;
    if (arc_index == 953) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 958) return "E"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 961) return "E"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 965) return "E"  ;
    if (arc_index == 967) return "E"  ;
    if (arc_index == 1013) return "H"  ;
    if (arc_index == 1018) return "H"  ;
    if (arc_index == 1056) return "H"  ;
    if (arc_index == 1078) return "E"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1081) return "E"  ;
    if (arc_index == 1082) return "E"  ;
    if (arc_index == 1083) return "E"  ;
    if (arc_index == 1084) return "E"  ;
    if (arc_index == 1085) return "E"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1087) return "E"  ;
    if (arc_index == 1088) return "E"  ;
    if (arc_index == 1089) return "E"  ;
    if (arc_index == 1090) return "E"  ;
    if (arc_index == 1091) return "E"  ;
    if (arc_index == 1092) return "E"  ;
    if (arc_index == 1093) return "E"  ;
    if (arc_index == 1094) return "E"  ;
    if (arc_index == 1095) return "E"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1097) return "E"  ;
    if (arc_index == 1098) return "E"  ;
    if (arc_index == 1099) return "E"  ;
    if (arc_index == 1111) return "H"  ;
    if (arc_index == 1156) return "H"  ;
    if (arc_index == 1224) return "E"  ;
    if (arc_index == 1355) return "H"  ;
    if (arc_index == 1400) return "W"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1484) return "W"  ;
    if (arc_index == 1532) return "H"  ;
    if (arc_index == 1600) return "H"  ;
    if (arc_index == 1601) return "H"  ;
    if (arc_index == 1616) return "H"  ;
    if (arc_index == 1709) return "W"  ;
    if (arc_index == 1722) return "W"  ;
    if (arc_index == 1725) return "H"  ;
    if (arc_index == 1733) return "W"  ;
    if (arc_index == 1748) return "W"  ;
    if (arc_index == 1798) return "W"  ;
    if (arc_index == 1808) return "W"  ;
    if (arc_index == 1812) return "W"  ;
    if (arc_index == 1841) return "H"  ;
    if (arc_index == 1889) return "H"  ;
    if (arc_index == 1897) return "H"  ;
    if (arc_index == 1930) return "H"  ;
    if (arc_index == 1934) return "H"  ;
    if (arc_index == 1944) return "H"  ;
    if (arc_index == 1955) return "H"  ;
    if (arc_index == 1957) return "H"  ;
    if (arc_index == 2038) return "H"  ;
    if (arc_index == 2075) return "H"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2115) return "W"  ;
    if (arc_index == 2176) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2228) return "H"  ;
    if (arc_index == 2232) return "H"  ;
    if (arc_index == 2305) return "H"  ;
    if (arc_index == 2474) return "H"  ;
    if (arc_index == 2552) return "H"  ;
    if (arc_index == 2555) return "H"  ;
    if (arc_index == 2556) return "H"  ;
    if (arc_index == 2557) return "E"  ;
    if (arc_index == 2561) return "E"  ;
    if (arc_index == 2566) return "E"  ;
    if (arc_index == 2571) return "E"  ;
    if (arc_index == 2585) return "E"  ;
    if (arc_index == 2730) return "E"  ;
    if (arc_index == 2733) return "E"  ;
    if (arc_index == 2734) return "W"  ;
    if (arc_index == 2740) return "W"  ;
    if (arc_index == 2746) return "W"  ;
    if (arc_index == 2747) return "W"  ;
    if (arc_index == 2748) return "W"  ;
    if (arc_index == 2761) return "W"  ;
    if (arc_index == 2792) return "W"  ;
    if (arc_index == 2796) return "W"  ;
    if (arc_index == 2800) return "E"  ;
    if (arc_index == 2802) return "E"  ;
    if (arc_index == 2803) return "E"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2809) return "E"  ;
    if (arc_index == 2811) return "E"  ;
    if (arc_index == 2812) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2814) return "E"  ;
    if (arc_index == 2851) return "E"  ;
    if (arc_index == 2859) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2877) return "H"  ;
    if (arc_index == 2900) return "W"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 6)) begin 
    if (arc_index == 4) return "W"  ;
    if (arc_index == 5) return "W"  ;
    if (arc_index == 6) return "W"  ;
    if (arc_index == 9) return "W"  ;
    if (arc_index == 12) return "W"  ;
    if (arc_index == 14) return "W"  ;
    if (arc_index == 16) return "W"  ;
    if (arc_index == 28) return "E"  ;
    if (arc_index == 30) return "E"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 113) return "E"  ;
    if (arc_index == 125) return "E"  ;
    if (arc_index == 128) return "H"  ;
    if (arc_index == 158) return "H"  ;
    if (arc_index == 159) return "H"  ;
    if (arc_index == 160) return "H"  ;
    if (arc_index == 205) return "H"  ;
    if (arc_index == 210) return "H"  ;
    if (arc_index == 212) return "H"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 261) return "H"  ;
    if (arc_index == 269) return "H"  ;
    if (arc_index == 273) return "H"  ;
    if (arc_index == 278) return "H"  ;
    if (arc_index == 327) return "H"  ;
    if (arc_index == 340) return "H"  ;
    if (arc_index == 356) return "H"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 399) return "E"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 426) return "E"  ;
    if (arc_index == 436) return "E"  ;
    if (arc_index == 482) return "H"  ;
    if (arc_index == 485) return "H"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 593) return "H"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 642) return "W"  ;
    if (arc_index == 649) return "E"  ;
    if (arc_index == 655) return "E"  ;
    if (arc_index == 663) return "H"  ;
    if (arc_index == 686) return "H"  ;
    if (arc_index == 691) return "H"  ;
    if (arc_index == 706) return "H"  ;
    if (arc_index == 721) return "W"  ;
    if (arc_index == 763) return "W"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 819) return "W"  ;
    if (arc_index == 822) return "W"  ;
    if (arc_index == 836) return "W"  ;
    if (arc_index == 837) return "W"  ;
    if (arc_index == 838) return "H"  ;
    if (arc_index == 839) return "H"  ;
    if (arc_index == 850) return "H"  ;
    if (arc_index == 851) return "H"  ;
    if (arc_index == 852) return "H"  ;
    if (arc_index == 857) return "E"  ;
    if (arc_index == 863) return "E"  ;
    if (arc_index == 869) return "E"  ;
    if (arc_index == 882) return "E"  ;
    if (arc_index == 883) return "E"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 965) return "E"  ;
    if (arc_index == 971) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1035) return "H"  ;
    if (arc_index == 1038) return "H"  ;
    if (arc_index == 1056) return "W"  ;
    if (arc_index == 1062) return "W"  ;
    if (arc_index == 1078) return "H"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1089) return "E"  ;
    if (arc_index == 1100) return "E"  ;
    if (arc_index == 1101) return "E"  ;
    if (arc_index == 1102) return "E"  ;
    if (arc_index == 1103) return "E"  ;
    if (arc_index == 1104) return "W"  ;
    if (arc_index == 1105) return "W"  ;
    if (arc_index == 1106) return "W"  ;
    if (arc_index == 1107) return "W"  ;
    if (arc_index == 1108) return "W"  ;
    if (arc_index == 1109) return "W"  ;
    if (arc_index == 1110) return "W"  ;
    if (arc_index == 1111) return "W"  ;
    if (arc_index == 1112) return "W"  ;
    if (arc_index == 1113) return "W"  ;
    if (arc_index == 1114) return "W"  ;
    if (arc_index == 1115) return "W"  ;
    if (arc_index == 1116) return "W"  ;
    if (arc_index == 1117) return "W"  ;
    if (arc_index == 1118) return "E"  ;
    if (arc_index == 1119) return "E"  ;
    if (arc_index == 1120) return "E"  ;
    if (arc_index == 1121) return "W"  ;
    if (arc_index == 1124) return "W"  ;
    if (arc_index == 1133) return "H"  ;
    if (arc_index == 1149) return "W"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1164) return "W"  ;
    if (arc_index == 1174) return "W"  ;
    if (arc_index == 1178) return "H"  ;
    if (arc_index == 1187) return "H"  ;
    if (arc_index == 1190) return "H"  ;
    if (arc_index == 1195) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1275) return "E"  ;
    if (arc_index == 1286) return "E"  ;
    if (arc_index == 1290) return "E"  ;
    if (arc_index == 1334) return "E"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1341) return "W"  ;
    if (arc_index == 1344) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1377) return "H"  ;
    if (arc_index == 1394) return "E"  ;
    if (arc_index == 1396) return "E"  ;
    if (arc_index == 1398) return "E"  ;
    if (arc_index == 1401) return "E"  ;
    if (arc_index == 1405) return "E"  ;
    if (arc_index == 1413) return "E"  ;
    if (arc_index == 1415) return "E"  ;
    if (arc_index == 1422) return "E"  ;
    if (arc_index == 1423) return "E"  ;
    if (arc_index == 1449) return "E"  ;
    if (arc_index == 1456) return "E"  ;
    if (arc_index == 1462) return "E"  ;
    if (arc_index == 1470) return "E"  ;
    if (arc_index == 1471) return "E"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1541) return "W"  ;
    if (arc_index == 1543) return "W"  ;
    if (arc_index == 1554) return "H"  ;
    if (arc_index == 1580) return "H"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1610) return "E"  ;
    if (arc_index == 1613) return "E"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1619) return "E"  ;
    if (arc_index == 1620) return "E"  ;
    if (arc_index == 1638) return "H"  ;
    if (arc_index == 1650) return "H"  ;
    if (arc_index == 1653) return "E"  ;
    if (arc_index == 1654) return "E"  ;
    if (arc_index == 1691) return "W"  ;
    if (arc_index == 1703) return "W"  ;
    if (arc_index == 1704) return "W"  ;
    if (arc_index == 1736) return "E"  ;
    if (arc_index == 1737) return "E"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1747) return "H"  ;
    if (arc_index == 1773) return "W"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1782) return "E"  ;
    if (arc_index == 1785) return "E"  ;
    if (arc_index == 1787) return "E"  ;
    if (arc_index == 1788) return "E"  ;
    if (arc_index == 1789) return "W"  ;
    if (arc_index == 1790) return "W"  ;
    if (arc_index == 1792) return "E"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1799) return "W"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1802) return "W"  ;
    if (arc_index == 1803) return "E"  ;
    if (arc_index == 1804) return "W"  ;
    if (arc_index == 1808) return "W"  ;
    if (arc_index == 1812) return "W"  ;
    if (arc_index == 1815) return "W"  ;
    if (arc_index == 1822) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1829) return "W"  ;
    if (arc_index == 1847) return "E"  ;
    if (arc_index == 1848) return "E"  ;
    if (arc_index == 1851) return "E"  ;
    if (arc_index == 1858) return "E"  ;
    if (arc_index == 1860) return "E"  ;
    if (arc_index == 1863) return "H"  ;
    if (arc_index == 1867) return "E"  ;
    if (arc_index == 1869) return "E"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1906) return "W"  ;
    if (arc_index == 1917) return "E"  ;
    if (arc_index == 1928) return "E"  ;
    if (arc_index == 1952) return "H"  ;
    if (arc_index == 1966) return "H"  ;
    if (arc_index == 1979) return "H"  ;
    if (arc_index == 1988) return "H"  ;
    if (arc_index == 1994) return "H"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2059) return "E"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2090) return "W"  ;
    if (arc_index == 2091) return "W"  ;
    if (arc_index == 2095) return "W"  ;
    if (arc_index == 2097) return "H"  ;
    if (arc_index == 2121) return "E"  ;
    if (arc_index == 2152) return "E"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2237) return "E"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2250) return "H"  ;
    if (arc_index == 2252) return "H"  ;
    if (arc_index == 2257) return "W"  ;
    if (arc_index == 2260) return "W"  ;
    if (arc_index == 2262) return "W"  ;
    if (arc_index == 2265) return "W"  ;
    if (arc_index == 2268) return "W"  ;
    if (arc_index == 2274) return "W"  ;
    if (arc_index == 2280) return "W"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2302) return "W"  ;
    if (arc_index == 2308) return "W"  ;
    if (arc_index == 2313) return "W"  ;
    if (arc_index == 2318) return "W"  ;
    if (arc_index == 2320) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2346) return "W"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2363) return "W"  ;
    if (arc_index == 2368) return "W"  ;
    if (arc_index == 2369) return "W"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2375) return "W"  ;
    if (arc_index == 2386) return "W"  ;
    if (arc_index == 2413) return "W"  ;
    if (arc_index == 2424) return "E"  ;
    if (arc_index == 2429) return "E"  ;
    if (arc_index == 2449) return "E"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2507) return "E"  ;
    if (arc_index == 2543) return "E"  ;
    if (arc_index == 2548) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2611) return "W"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2627) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2687) return "W"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2714) return "W"  ;
    if (arc_index == 2738) return "W"  ;
    if (arc_index == 2749) return "W"  ;
    if (arc_index == 2782) return "W"  ;
    if (arc_index == 2784) return "W"  ;
    if (arc_index == 2801) return "E"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2817) return "W"  ;
    if (arc_index == 2840) return "W"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2892) return "E"  ;
    if (arc_index == 2894) return "E"  ;
    if (arc_index == 2899) return "H"  ;
    if (arc_index == 2919) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 10)) begin 
    if (arc_index == 146) return "W"  ;
    if (arc_index == 150) return "H"  ;
    if (arc_index == 283) return "H"  ;
    if (arc_index == 289) return "W"  ;
    if (arc_index == 291) return "H"  ;
    if (arc_index == 378) return "H"  ;
    if (arc_index == 416) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 504) return "H"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 615) return "H"  ;
    if (arc_index == 685) return "H"  ;
    if (arc_index == 723) return "H"  ;
    if (arc_index == 818) return "H"  ;
    if (arc_index == 860) return "H"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1035) return "W"  ;
    if (arc_index == 1036) return "W"  ;
    if (arc_index == 1039) return "W"  ;
    if (arc_index == 1040) return "W"  ;
    if (arc_index == 1041) return "W"  ;
    if (arc_index == 1043) return "W"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1046) return "W"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1055) return "W"  ;
    if (arc_index == 1057) return "H"  ;
    if (arc_index == 1100) return "H"  ;
    if (arc_index == 1122) return "H"  ;
    if (arc_index == 1123) return "W"  ;
    if (arc_index == 1124) return "W"  ;
    if (arc_index == 1125) return "W"  ;
    if (arc_index == 1126) return "W"  ;
    if (arc_index == 1127) return "W"  ;
    if (arc_index == 1128) return "W"  ;
    if (arc_index == 1129) return "W"  ;
    if (arc_index == 1130) return "W"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1132) return "W"  ;
    if (arc_index == 1133) return "W"  ;
    if (arc_index == 1134) return "W"  ;
    if (arc_index == 1135) return "W"  ;
    if (arc_index == 1136) return "W"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1138) return "W"  ;
    if (arc_index == 1139) return "W"  ;
    if (arc_index == 1140) return "W"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1142) return "W"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1155) return "H"  ;
    if (arc_index == 1200) return "H"  ;
    if (arc_index == 1300) return "H"  ;
    if (arc_index == 1311) return "E"  ;
    if (arc_index == 1399) return "H"  ;
    if (arc_index == 1540) return "H"  ;
    if (arc_index == 1566) return "W"  ;
    if (arc_index == 1567) return "W"  ;
    if (arc_index == 1570) return "W"  ;
    if (arc_index == 1572) return "E"  ;
    if (arc_index == 1573) return "E"  ;
    if (arc_index == 1575) return "W"  ;
    if (arc_index == 1576) return "H"  ;
    if (arc_index == 1577) return "H"  ;
    if (arc_index == 1579) return "H"  ;
    if (arc_index == 1580) return "H"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1582) return "W"  ;
    if (arc_index == 1583) return "W"  ;
    if (arc_index == 1595) return "W"  ;
    if (arc_index == 1660) return "H"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1769) return "H"  ;
    if (arc_index == 1839) return "H"  ;
    if (arc_index == 1885) return "H"  ;
    if (arc_index == 1900) return "E"  ;
    if (arc_index == 1974) return "H"  ;
    if (arc_index == 1988) return "H"  ;
    if (arc_index == 2003) return "H"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2100) return "W"  ;
    if (arc_index == 2119) return "H"  ;
    if (arc_index == 2178) return "W"  ;
    if (arc_index == 2184) return "E"  ;
    if (arc_index == 2203) return "E"  ;
    if (arc_index == 2211) return "E"  ;
    if (arc_index == 2272) return "H"  ;
    if (arc_index == 2414) return "H"  ;
    if (arc_index == 2559) return "H"  ;
    if (arc_index == 2595) return "H"  ;
    if (arc_index == 2650) return "H"  ;
    if (arc_index == 2654) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2712) return "W"  ;
    if (arc_index == 2726) return "W"  ;
    if (arc_index == 2921) return "H"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 10)) begin 
    if (arc_index == 17) return "H"  ;
    if (arc_index == 46) return "H"  ;
    if (arc_index == 172) return "H"  ;
    if (arc_index == 179) return "E"  ;
    if (arc_index == 191) return "W"  ;
    if (arc_index == 197) return "W"  ;
    if (arc_index == 203) return "W"  ;
    if (arc_index == 213) return "W"  ;
    if (arc_index == 254) return "W"  ;
    if (arc_index == 286) return "W"  ;
    if (arc_index == 288) return "W"  ;
    if (arc_index == 294) return "W"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 305) return "H"  ;
    if (arc_index == 307) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 313) return "H"  ;
    if (arc_index == 316) return "H"  ;
    if (arc_index == 318) return "E"  ;
    if (arc_index == 319) return "E"  ;
    if (arc_index == 324) return "E"  ;
    if (arc_index == 339) return "E"  ;
    if (arc_index == 341) return "E"  ;
    if (arc_index == 370) return "E"  ;
    if (arc_index == 400) return "H"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 526) return "H"  ;
    if (arc_index == 563) return "H"  ;
    if (arc_index == 568) return "E"  ;
    if (arc_index == 594) return "E"  ;
    if (arc_index == 598) return "E"  ;
    if (arc_index == 601) return "E"  ;
    if (arc_index == 616) return "E"  ;
    if (arc_index == 620) return "E"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 627) return "W"  ;
    if (arc_index == 636) return "W"  ;
    if (arc_index == 637) return "H"  ;
    if (arc_index == 639) return "H"  ;
    if (arc_index == 689) return "E"  ;
    if (arc_index == 704) return "E"  ;
    if (arc_index == 707) return "H"  ;
    if (arc_index == 714) return "H"  ;
    if (arc_index == 718) return "W"  ;
    if (arc_index == 723) return "W"  ;
    if (arc_index == 725) return "W"  ;
    if (arc_index == 737) return "W"  ;
    if (arc_index == 741) return "E"  ;
    if (arc_index == 824) return "E"  ;
    if (arc_index == 842) return "E"  ;
    if (arc_index == 882) return "H"  ;
    if (arc_index == 1050) return "W"  ;
    if (arc_index == 1071) return "W"  ;
    if (arc_index == 1079) return "H"  ;
    if (arc_index == 1103) return "E"  ;
    if (arc_index == 1122) return "H"  ;
    if (arc_index == 1141) return "H"  ;
    if (arc_index == 1144) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1146) return "W"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1148) return "W"  ;
    if (arc_index == 1149) return "W"  ;
    if (arc_index == 1150) return "W"  ;
    if (arc_index == 1151) return "W"  ;
    if (arc_index == 1152) return "W"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1154) return "W"  ;
    if (arc_index == 1155) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1158) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1160) return "W"  ;
    if (arc_index == 1161) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1164) return "W"  ;
    if (arc_index == 1165) return "W"  ;
    if (arc_index == 1177) return "H"  ;
    if (arc_index == 1222) return "H"  ;
    if (arc_index == 1242) return "H"  ;
    if (arc_index == 1277) return "H"  ;
    if (arc_index == 1305) return "H"  ;
    if (arc_index == 1320) return "H"  ;
    if (arc_index == 1342) return "H"  ;
    if (arc_index == 1347) return "H"  ;
    if (arc_index == 1354) return "H"  ;
    if (arc_index == 1357) return "H"  ;
    if (arc_index == 1361) return "H"  ;
    if (arc_index == 1421) return "H"  ;
    if (arc_index == 1552) return "H"  ;
    if (arc_index == 1558) return "W"  ;
    if (arc_index == 1570) return "W"  ;
    if (arc_index == 1598) return "H"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1682) return "H"  ;
    if (arc_index == 1787) return "E"  ;
    if (arc_index == 1791) return "H"  ;
    if (arc_index == 1817) return "E"  ;
    if (arc_index == 1907) return "H"  ;
    if (arc_index == 1996) return "H"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2010) return "H"  ;
    if (arc_index == 2089) return "W"  ;
    if (arc_index == 2101) return "W"  ;
    if (arc_index == 2141) return "H"  ;
    if (arc_index == 2181) return "E"  ;
    if (arc_index == 2192) return "E"  ;
    if (arc_index == 2194) return "E"  ;
    if (arc_index == 2196) return "E"  ;
    if (arc_index == 2198) return "E"  ;
    if (arc_index == 2208) return "E"  ;
    if (arc_index == 2294) return "H"  ;
    if (arc_index == 2354) return "H"  ;
    if (arc_index == 2356) return "E"  ;
    if (arc_index == 2373) return "E"  ;
    if (arc_index == 2387) return "W"  ;
    if (arc_index == 2395) return "W"  ;
    if (arc_index == 2403) return "W"  ;
    if (arc_index == 2415) return "E"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2620) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2624) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2627) return "W"  ;
    if (arc_index == 2631) return "W"  ;
    if (arc_index == 2634) return "W"  ;
    if (arc_index == 2696) return "E"  ;
    if (arc_index == 2727) return "E"  ;
    if (arc_index == 2833) return "E"  ;
    if (arc_index == 2895) return "E"  ;
    if (arc_index == 2922) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 6)) begin 
    if (arc_index == 19) return "W"  ;
    if (arc_index == 20) return "W"  ;
    if (arc_index == 24) return "E"  ;
    if (arc_index == 29) return "E"  ;
    if (arc_index == 31) return "E"  ;
    if (arc_index == 39) return "H"  ;
    if (arc_index == 98) return "H"  ;
    if (arc_index == 100) return "W"  ;
    if (arc_index == 106) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 113) return "W"  ;
    if (arc_index == 118) return "E"  ;
    if (arc_index == 119) return "E"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 149) return "E"  ;
    if (arc_index == 163) return "W"  ;
    if (arc_index == 165) return "W"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 180) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 188) return "W"  ;
    if (arc_index == 194) return "H"  ;
    if (arc_index == 201) return "H"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 223) return "W"  ;
    if (arc_index == 224) return "W"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 229) return "W"  ;
    if (arc_index == 279) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 299) return "W"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 327) return "H"  ;
    if (arc_index == 330) return "H"  ;
    if (arc_index == 331) return "H"  ;
    if (arc_index == 335) return "H"  ;
    if (arc_index == 345) return "W"  ;
    if (arc_index == 351) return "W"  ;
    if (arc_index == 356) return "W"  ;
    if (arc_index == 359) return "E"  ;
    if (arc_index == 362) return "W"  ;
    if (arc_index == 363) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 367) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 402) return "E"  ;
    if (arc_index == 408) return "E"  ;
    if (arc_index == 422) return "H"  ;
    if (arc_index == 426) return "H"  ;
    if (arc_index == 436) return "H"  ;
    if (arc_index == 445) return "E"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 531) return "W"  ;
    if (arc_index == 548) return "H"  ;
    if (arc_index == 564) return "H"  ;
    if (arc_index == 595) return "H"  ;
    if (arc_index == 629) return "H"  ;
    if (arc_index == 639) return "H"  ;
    if (arc_index == 642) return "H"  ;
    if (arc_index == 647) return "H"  ;
    if (arc_index == 649) return "H"  ;
    if (arc_index == 653) return "H"  ;
    if (arc_index == 654) return "H"  ;
    if (arc_index == 655) return "H"  ;
    if (arc_index == 656) return "H"  ;
    if (arc_index == 658) return "E"  ;
    if (arc_index == 659) return "H"  ;
    if (arc_index == 660) return "E"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 677) return "E"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 726) return "W"  ;
    if (arc_index == 729) return "H"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 759) return "E"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 836) return "W"  ;
    if (arc_index == 850) return "W"  ;
    if (arc_index == 863) return "W"  ;
    if (arc_index == 866) return "W"  ;
    if (arc_index == 868) return "W"  ;
    if (arc_index == 869) return "W"  ;
    if (arc_index == 876) return "W"  ;
    if (arc_index == 890) return "W"  ;
    if (arc_index == 898) return "E"  ;
    if (arc_index == 904) return "H"  ;
    if (arc_index == 930) return "H"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 969) return "E"  ;
    if (arc_index == 977) return "E"  ;
    if (arc_index == 982) return "E"  ;
    if (arc_index == 997) return "E"  ;
    if (arc_index == 1014) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1044) return "E"  ;
    if (arc_index == 1046) return "W"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1059) return "W"  ;
    if (arc_index == 1069) return "W"  ;
    if (arc_index == 1085) return "W"  ;
    if (arc_index == 1092) return "W"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1100) return "E"  ;
    if (arc_index == 1101) return "H"  ;
    if (arc_index == 1102) return "H"  ;
    if (arc_index == 1107) return "H"  ;
    if (arc_index == 1114) return "H"  ;
    if (arc_index == 1115) return "H"  ;
    if (arc_index == 1144) return "H"  ;
    if (arc_index == 1162) return "H"  ;
    if (arc_index == 1166) return "W"  ;
    if (arc_index == 1167) return "E"  ;
    if (arc_index == 1168) return "E"  ;
    if (arc_index == 1169) return "W"  ;
    if (arc_index == 1170) return "W"  ;
    if (arc_index == 1171) return "W"  ;
    if (arc_index == 1172) return "W"  ;
    if (arc_index == 1173) return "E"  ;
    if (arc_index == 1174) return "E"  ;
    if (arc_index == 1175) return "E"  ;
    if (arc_index == 1176) return "E"  ;
    if (arc_index == 1177) return "E"  ;
    if (arc_index == 1178) return "E"  ;
    if (arc_index == 1179) return "W"  ;
    if (arc_index == 1180) return "W"  ;
    if (arc_index == 1181) return "W"  ;
    if (arc_index == 1182) return "W"  ;
    if (arc_index == 1183) return "E"  ;
    if (arc_index == 1184) return "W"  ;
    if (arc_index == 1185) return "W"  ;
    if (arc_index == 1186) return "W"  ;
    if (arc_index == 1187) return "W"  ;
    if (arc_index == 1189) return "W"  ;
    if (arc_index == 1199) return "H"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1211) return "E"  ;
    if (arc_index == 1217) return "E"  ;
    if (arc_index == 1218) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1244) return "H"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1266) return "W"  ;
    if (arc_index == 1272) return "W"  ;
    if (arc_index == 1279) return "W"  ;
    if (arc_index == 1288) return "W"  ;
    if (arc_index == 1289) return "W"  ;
    if (arc_index == 1292) return "W"  ;
    if (arc_index == 1293) return "W"  ;
    if (arc_index == 1295) return "W"  ;
    if (arc_index == 1296) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1365) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1368) return "W"  ;
    if (arc_index == 1377) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1396) return "W"  ;
    if (arc_index == 1401) return "W"  ;
    if (arc_index == 1433) return "E"  ;
    if (arc_index == 1442) return "E"  ;
    if (arc_index == 1443) return "H"  ;
    if (arc_index == 1456) return "H"  ;
    if (arc_index == 1471) return "E"  ;
    if (arc_index == 1474) return "E"  ;
    if (arc_index == 1490) return "E"  ;
    if (arc_index == 1500) return "E"  ;
    if (arc_index == 1507) return "E"  ;
    if (arc_index == 1515) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1546) return "W"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1620) return "H"  ;
    if (arc_index == 1631) return "H"  ;
    if (arc_index == 1640) return "H"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1687) return "E"  ;
    if (arc_index == 1704) return "H"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1764) return "E"  ;
    if (arc_index == 1788) return "E"  ;
    if (arc_index == 1813) return "H"  ;
    if (arc_index == 1820) return "W"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1871) return "E"  ;
    if (arc_index == 1872) return "W"  ;
    if (arc_index == 1878) return "W"  ;
    if (arc_index == 1881) return "W"  ;
    if (arc_index == 1883) return "W"  ;
    if (arc_index == 1884) return "W"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 1923) return "E"  ;
    if (arc_index == 1929) return "H"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1965) return "W"  ;
    if (arc_index == 1976) return "W"  ;
    if (arc_index == 1988) return "E"  ;
    if (arc_index == 2018) return "H"  ;
    if (arc_index == 2032) return "H"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2120) return "W"  ;
    if (arc_index == 2127) return "W"  ;
    if (arc_index == 2130) return "E"  ;
    if (arc_index == 2133) return "E"  ;
    if (arc_index == 2141) return "E"  ;
    if (arc_index == 2163) return "H"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2246) return "E"  ;
    if (arc_index == 2251) return "E"  ;
    if (arc_index == 2306) return "E"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2316) return "H"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2330) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2398) return "W"  ;
    if (arc_index == 2426) return "E"  ;
    if (arc_index == 2428) return "E"  ;
    if (arc_index == 2431) return "E"  ;
    if (arc_index == 2435) return "E"  ;
    if (arc_index == 2439) return "E"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2505) return "E"  ;
    if (arc_index == 2512) return "E"  ;
    if (arc_index == 2521) return "E"  ;
    if (arc_index == 2524) return "E"  ;
    if (arc_index == 2528) return "E"  ;
    if (arc_index == 2534) return "E"  ;
    if (arc_index == 2599) return "E"  ;
    if (arc_index == 2614) return "E"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2736) return "E"  ;
    if (arc_index == 2752) return "E"  ;
    if (arc_index == 2771) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2820) return "E"  ;
    if (arc_index == 2841) return "E"  ;
    if (arc_index == 2922) return "W"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 2)) begin 
    if (arc_index == 61) return "H"  ;
    if (arc_index == 67) return "H"  ;
    if (arc_index == 73) return "H"  ;
    if (arc_index == 85) return "H"  ;
    if (arc_index == 99) return "H"  ;
    if (arc_index == 115) return "H"  ;
    if (arc_index == 144) return "H"  ;
    if (arc_index == 145) return "H"  ;
    if (arc_index == 216) return "H"  ;
    if (arc_index == 238) return "W"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 349) return "H"  ;
    if (arc_index == 357) return "H"  ;
    if (arc_index == 371) return "W"  ;
    if (arc_index == 444) return "H"  ;
    if (arc_index == 451) return "H"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 466) return "W"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 491) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 530) return "E"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 570) return "H"  ;
    if (arc_index == 640) return "H"  ;
    if (arc_index == 641) return "H"  ;
    if (arc_index == 679) return "W"  ;
    if (arc_index == 681) return "H"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 750) return "W"  ;
    if (arc_index == 751) return "H"  ;
    if (arc_index == 770) return "H"  ;
    if (arc_index == 779) return "E"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 797) return "E"  ;
    if (arc_index == 799) return "E"  ;
    if (arc_index == 800) return "W"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 803) return "E"  ;
    if (arc_index == 808) return "E"  ;
    if (arc_index == 809) return "E"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 811) return "E"  ;
    if (arc_index == 812) return "E"  ;
    if (arc_index == 865) return "E"  ;
    if (arc_index == 900) return "W"  ;
    if (arc_index == 902) return "W"  ;
    if (arc_index == 915) return "E"  ;
    if (arc_index == 924) return "E"  ;
    if (arc_index == 926) return "H"  ;
    if (arc_index == 928) return "E"  ;
    if (arc_index == 931) return "E"  ;
    if (arc_index == 932) return "E"  ;
    if (arc_index == 935) return "E"  ;
    if (arc_index == 938) return "E"  ;
    if (arc_index == 942) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 957) return "E"  ;
    if (arc_index == 978) return "E"  ;
    if (arc_index == 979) return "W"  ;
    if (arc_index == 1011) return "W"  ;
    if (arc_index == 1016) return "W"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1032) return "E"  ;
    if (arc_index == 1123) return "H"  ;
    if (arc_index == 1166) return "H"  ;
    if (arc_index == 1179) return "H"  ;
    if (arc_index == 1188) return "W"  ;
    if (arc_index == 1189) return "E"  ;
    if (arc_index == 1190) return "E"  ;
    if (arc_index == 1191) return "E"  ;
    if (arc_index == 1192) return "E"  ;
    if (arc_index == 1193) return "E"  ;
    if (arc_index == 1194) return "E"  ;
    if (arc_index == 1195) return "E"  ;
    if (arc_index == 1196) return "E"  ;
    if (arc_index == 1197) return "E"  ;
    if (arc_index == 1198) return "E"  ;
    if (arc_index == 1199) return "E"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1201) return "E"  ;
    if (arc_index == 1202) return "E"  ;
    if (arc_index == 1203) return "W"  ;
    if (arc_index == 1204) return "E"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1207) return "E"  ;
    if (arc_index == 1208) return "E"  ;
    if (arc_index == 1209) return "E"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1211) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1214) return "E"  ;
    if (arc_index == 1215) return "E"  ;
    if (arc_index == 1217) return "E"  ;
    if (arc_index == 1218) return "E"  ;
    if (arc_index == 1221) return "H"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1230) return "E"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1266) return "H"  ;
    if (arc_index == 1288) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1462) return "W"  ;
    if (arc_index == 1465) return "H"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1496) return "W"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1522) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1528) return "E"  ;
    if (arc_index == 1529) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1533) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1539) return "E"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1589) return "E"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1603) return "E"  ;
    if (arc_index == 1642) return "H"  ;
    if (arc_index == 1644) return "H"  ;
    if (arc_index == 1658) return "H"  ;
    if (arc_index == 1723) return "E"  ;
    if (arc_index == 1726) return "H"  ;
    if (arc_index == 1735) return "W"  ;
    if (arc_index == 1740) return "W"  ;
    if (arc_index == 1743) return "W"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1789) return "E"  ;
    if (arc_index == 1790) return "E"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1835) return "H"  ;
    if (arc_index == 1857) return "W"  ;
    if (arc_index == 1864) return "W"  ;
    if (arc_index == 1921) return "W"  ;
    if (arc_index == 1935) return "W"  ;
    if (arc_index == 1937) return "W"  ;
    if (arc_index == 1951) return "H"  ;
    if (arc_index == 1972) return "W"  ;
    if (arc_index == 1973) return "W"  ;
    if (arc_index == 2002) return "W"  ;
    if (arc_index == 2006) return "E"  ;
    if (arc_index == 2007) return "E"  ;
    if (arc_index == 2013) return "E"  ;
    if (arc_index == 2014) return "E"  ;
    if (arc_index == 2015) return "E"  ;
    if (arc_index == 2020) return "E"  ;
    if (arc_index == 2021) return "E"  ;
    if (arc_index == 2023) return "E"  ;
    if (arc_index == 2035) return "E"  ;
    if (arc_index == 2040) return "H"  ;
    if (arc_index == 2054) return "H"  ;
    if (arc_index == 2056) return "W"  ;
    if (arc_index == 2062) return "W"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2162) return "W"  ;
    if (arc_index == 2185) return "H"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2281) return "W"  ;
    if (arc_index == 2338) return "H"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2436) return "W"  ;
    if (arc_index == 2452) return "W"  ;
    if (arc_index == 2526) return "W"  ;
    if (arc_index == 2527) return "W"  ;
    if (arc_index == 2584) return "E"  ;
    if (arc_index == 2589) return "E"  ;
    if (arc_index == 2640) return "E"  ;
    if (arc_index == 2672) return "E"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2723) return "E"  ;
    if (arc_index == 2733) return "E"  ;
    if (arc_index == 2746) return "E"  ;
    if (arc_index == 2747) return "E"  ;
    if (arc_index == 2765) return "E"  ;
    if (arc_index == 2793) return "W"  ;
    if (arc_index == 2868) return "W"  ;
    if (arc_index == 2874) return "E"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2887) return "E"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 1)) begin 
    if (arc_index == 83) return "H"  ;
    if (arc_index == 135) return "W"  ;
    if (arc_index == 238) return "H"  ;
    if (arc_index == 268) return "H"  ;
    if (arc_index == 309) return "H"  ;
    if (arc_index == 371) return "H"  ;
    if (arc_index == 375) return "H"  ;
    if (arc_index == 379) return "H"  ;
    if (arc_index == 380) return "H"  ;
    if (arc_index == 384) return "H"  ;
    if (arc_index == 388) return "H"  ;
    if (arc_index == 389) return "H"  ;
    if (arc_index == 390) return "H"  ;
    if (arc_index == 391) return "W"  ;
    if (arc_index == 395) return "W"  ;
    if (arc_index == 418) return "W"  ;
    if (arc_index == 451) return "E"  ;
    if (arc_index == 452) return "E"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 466) return "H"  ;
    if (arc_index == 487) return "H"  ;
    if (arc_index == 491) return "E"  ;
    if (arc_index == 513) return "E"  ;
    if (arc_index == 514) return "E"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 575) return "W"  ;
    if (arc_index == 592) return "H"  ;
    if (arc_index == 679) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 703) return "H"  ;
    if (arc_index == 750) return "H"  ;
    if (arc_index == 773) return "H"  ;
    if (arc_index == 800) return "H"  ;
    if (arc_index == 900) return "W"  ;
    if (arc_index == 912) return "W"  ;
    if (arc_index == 948) return "H"  ;
    if (arc_index == 979) return "H"  ;
    if (arc_index == 1011) return "W"  ;
    if (arc_index == 1013) return "W"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1017) return "E"  ;
    if (arc_index == 1018) return "E"  ;
    if (arc_index == 1024) return "E"  ;
    if (arc_index == 1026) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1029) return "E"  ;
    if (arc_index == 1090) return "E"  ;
    if (arc_index == 1145) return "H"  ;
    if (arc_index == 1188) return "H"  ;
    if (arc_index == 1203) return "H"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1211) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1213) return "E"  ;
    if (arc_index == 1214) return "E"  ;
    if (arc_index == 1215) return "E"  ;
    if (arc_index == 1216) return "E"  ;
    if (arc_index == 1217) return "E"  ;
    if (arc_index == 1218) return "E"  ;
    if (arc_index == 1219) return "E"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1221) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1223) return "E"  ;
    if (arc_index == 1224) return "E"  ;
    if (arc_index == 1225) return "E"  ;
    if (arc_index == 1226) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1230) return "E"  ;
    if (arc_index == 1231) return "E"  ;
    if (arc_index == 1243) return "H"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1288) return "H"  ;
    if (arc_index == 1372) return "H"  ;
    if (arc_index == 1466) return "H"  ;
    if (arc_index == 1487) return "H"  ;
    if (arc_index == 1496) return "W"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1522) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1524) return "E"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1528) return "E"  ;
    if (arc_index == 1529) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1533) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1539) return "E"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1589) return "E"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1602) return "E"  ;
    if (arc_index == 1603) return "E"  ;
    if (arc_index == 1659) return "E"  ;
    if (arc_index == 1664) return "H"  ;
    if (arc_index == 1735) return "H"  ;
    if (arc_index == 1748) return "H"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1830) return "W"  ;
    if (arc_index == 1857) return "H"  ;
    if (arc_index == 1942) return "H"  ;
    if (arc_index == 1951) return "E"  ;
    if (arc_index == 1956) return "E"  ;
    if (arc_index == 1972) return "W"  ;
    if (arc_index == 1973) return "H"  ;
    if (arc_index == 2056) return "W"  ;
    if (arc_index == 2062) return "H"  ;
    if (arc_index == 2076) return "H"  ;
    if (arc_index == 2173) return "H"  ;
    if (arc_index == 2207) return "H"  ;
    if (arc_index == 2230) return "H"  ;
    if (arc_index == 2281) return "W"  ;
    if (arc_index == 2360) return "H"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2436) return "W"  ;
    if (arc_index == 2469) return "W"  ;
    if (arc_index == 2552) return "W"  ;
    if (arc_index == 2556) return "W"  ;
    if (arc_index == 2574) return "W"  ;
    if (arc_index == 2576) return "W"  ;
    if (arc_index == 2579) return "W"  ;
    if (arc_index == 2580) return "W"  ;
    if (arc_index == 2582) return "W"  ;
    if (arc_index == 2583) return "W"  ;
    if (arc_index == 2585) return "W"  ;
    if (arc_index == 2589) return "E"  ;
    if (arc_index == 2590) return "E"  ;
    if (arc_index == 2593) return "E"  ;
    if (arc_index == 2607) return "E"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2682) return "E"  ;
    if (arc_index == 2747) return "E"  ;
    if (arc_index == 2793) return "E"  ;
    if (arc_index == 2811) return "E"  ;
    if (arc_index == 2851) return "E"  ;
    if (arc_index == 2863) return "E"  ;
    if (arc_index == 2874) return "E"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2879) return "E"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 9)) begin 
    if (arc_index == 8) return "E"  ;
    if (arc_index == 105) return "H"  ;
    if (arc_index == 139) return "E"  ;
    if (arc_index == 147) return "E"  ;
    if (arc_index == 171) return "E"  ;
    if (arc_index == 260) return "H"  ;
    if (arc_index == 326) return "H"  ;
    if (arc_index == 370) return "E"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 393) return "H"  ;
    if (arc_index == 401) return "H"  ;
    if (arc_index == 425) return "H"  ;
    if (arc_index == 427) return "E"  ;
    if (arc_index == 432) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 488) return "H"  ;
    if (arc_index == 527) return "H"  ;
    if (arc_index == 554) return "H"  ;
    if (arc_index == 614) return "H"  ;
    if (arc_index == 620) return "H"  ;
    if (arc_index == 672) return "H"  ;
    if (arc_index == 725) return "H"  ;
    if (arc_index == 740) return "E"  ;
    if (arc_index == 741) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 795) return "H"  ;
    if (arc_index == 871) return "H"  ;
    if (arc_index == 941) return "E"  ;
    if (arc_index == 970) return "H"  ;
    if (arc_index == 1035) return "H"  ;
    if (arc_index == 1039) return "W"  ;
    if (arc_index == 1040) return "W"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1126) return "W"  ;
    if (arc_index == 1167) return "H"  ;
    if (arc_index == 1200) return "H"  ;
    if (arc_index == 1210) return "H"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1232) return "W"  ;
    if (arc_index == 1233) return "W"  ;
    if (arc_index == 1234) return "W"  ;
    if (arc_index == 1235) return "W"  ;
    if (arc_index == 1236) return "W"  ;
    if (arc_index == 1237) return "E"  ;
    if (arc_index == 1238) return "W"  ;
    if (arc_index == 1239) return "W"  ;
    if (arc_index == 1240) return "W"  ;
    if (arc_index == 1241) return "E"  ;
    if (arc_index == 1242) return "E"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1244) return "W"  ;
    if (arc_index == 1245) return "W"  ;
    if (arc_index == 1246) return "W"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1248) return "W"  ;
    if (arc_index == 1249) return "E"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1251) return "W"  ;
    if (arc_index == 1252) return "W"  ;
    if (arc_index == 1253) return "W"  ;
    if (arc_index == 1265) return "H"  ;
    if (arc_index == 1298) return "H"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1302) return "W"  ;
    if (arc_index == 1303) return "W"  ;
    if (arc_index == 1304) return "W"  ;
    if (arc_index == 1305) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1309) return "W"  ;
    if (arc_index == 1310) return "H"  ;
    if (arc_index == 1313) return "H"  ;
    if (arc_index == 1316) return "H"  ;
    if (arc_index == 1331) return "H"  ;
    if (arc_index == 1342) return "H"  ;
    if (arc_index == 1509) return "H"  ;
    if (arc_index == 1566) return "H"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1686) return "H"  ;
    if (arc_index == 1752) return "H"  ;
    if (arc_index == 1770) return "H"  ;
    if (arc_index == 1836) return "H"  ;
    if (arc_index == 1879) return "H"  ;
    if (arc_index == 1900) return "H"  ;
    if (arc_index == 1974) return "H"  ;
    if (arc_index == 1995) return "H"  ;
    if (arc_index == 2046) return "E"  ;
    if (arc_index == 2069) return "W"  ;
    if (arc_index == 2071) return "W"  ;
    if (arc_index == 2074) return "W"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2084) return "H"  ;
    if (arc_index == 2086) return "W"  ;
    if (arc_index == 2098) return "H"  ;
    if (arc_index == 2146) return "E"  ;
    if (arc_index == 2180) return "E"  ;
    if (arc_index == 2195) return "W"  ;
    if (arc_index == 2197) return "W"  ;
    if (arc_index == 2208) return "E"  ;
    if (arc_index == 2229) return "H"  ;
    if (arc_index == 2272) return "H"  ;
    if (arc_index == 2295) return "H"  ;
    if (arc_index == 2325) return "H"  ;
    if (arc_index == 2377) return "H"  ;
    if (arc_index == 2382) return "H"  ;
    if (arc_index == 2396) return "W"  ;
    if (arc_index == 2455) return "W"  ;
    if (arc_index == 2522) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2655) return "W"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 8)) begin 
    if (arc_index == 89) return "W"  ;
    if (arc_index == 94) return "W"  ;
    if (arc_index == 104) return "W"  ;
    if (arc_index == 105) return "E"  ;
    if (arc_index == 111) return "E"  ;
    if (arc_index == 127) return "H"  ;
    if (arc_index == 147) return "E"  ;
    if (arc_index == 166) return "W"  ;
    if (arc_index == 171) return "E"  ;
    if (arc_index == 219) return "E"  ;
    if (arc_index == 240) return "E"  ;
    if (arc_index == 252) return "E"  ;
    if (arc_index == 260) return "E"  ;
    if (arc_index == 271) return "E"  ;
    if (arc_index == 282) return "H"  ;
    if (arc_index == 287) return "W"  ;
    if (arc_index == 364) return "W"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 393) return "E"  ;
    if (arc_index == 401) return "E"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 415) return "H"  ;
    if (arc_index == 423) return "H"  ;
    if (arc_index == 464) return "H"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 510) return "H"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 554) return "E"  ;
    if (arc_index == 596) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 636) return "H"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 704) return "E"  ;
    if (arc_index == 726) return "W"  ;
    if (arc_index == 729) return "W"  ;
    if (arc_index == 730) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 736) return "W"  ;
    if (arc_index == 737) return "W"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 740) return "E"  ;
    if (arc_index == 741) return "E"  ;
    if (arc_index == 742) return "W"  ;
    if (arc_index == 743) return "W"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 747) return "H"  ;
    if (arc_index == 759) return "H"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 795) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 817) return "H"  ;
    if (arc_index == 825) return "H"  ;
    if (arc_index == 867) return "H"  ;
    if (arc_index == 941) return "E"  ;
    if (arc_index == 970) return "E"  ;
    if (arc_index == 992) return "H"  ;
    if (arc_index == 1039) return "H"  ;
    if (arc_index == 1040) return "H"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1073) return "W"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1126) return "E"  ;
    if (arc_index == 1167) return "E"  ;
    if (arc_index == 1189) return "H"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1232) return "H"  ;
    if (arc_index == 1234) return "W"  ;
    if (arc_index == 1236) return "W"  ;
    if (arc_index == 1238) return "W"  ;
    if (arc_index == 1240) return "W"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1244) return "W"  ;
    if (arc_index == 1245) return "W"  ;
    if (arc_index == 1246) return "W"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1252) return "W"  ;
    if (arc_index == 1254) return "W"  ;
    if (arc_index == 1255) return "W"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1257) return "W"  ;
    if (arc_index == 1258) return "W"  ;
    if (arc_index == 1259) return "W"  ;
    if (arc_index == 1260) return "W"  ;
    if (arc_index == 1261) return "W"  ;
    if (arc_index == 1262) return "W"  ;
    if (arc_index == 1263) return "W"  ;
    if (arc_index == 1264) return "W"  ;
    if (arc_index == 1265) return "E"  ;
    if (arc_index == 1266) return "E"  ;
    if (arc_index == 1267) return "W"  ;
    if (arc_index == 1268) return "W"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1270) return "W"  ;
    if (arc_index == 1271) return "W"  ;
    if (arc_index == 1272) return "W"  ;
    if (arc_index == 1273) return "W"  ;
    if (arc_index == 1274) return "W"  ;
    if (arc_index == 1275) return "W"  ;
    if (arc_index == 1276) return "W"  ;
    if (arc_index == 1287) return "H"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1303) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1309) return "W"  ;
    if (arc_index == 1332) return "H"  ;
    if (arc_index == 1361) return "H"  ;
    if (arc_index == 1382) return "H"  ;
    if (arc_index == 1489) return "H"  ;
    if (arc_index == 1501) return "H"  ;
    if (arc_index == 1509) return "E"  ;
    if (arc_index == 1531) return "H"  ;
    if (arc_index == 1550) return "H"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1693) return "E"  ;
    if (arc_index == 1708) return "H"  ;
    if (arc_index == 1763) return "H"  ;
    if (arc_index == 1792) return "H"  ;
    if (arc_index == 1801) return "H"  ;
    if (arc_index == 1876) return "H"  ;
    if (arc_index == 1879) return "E"  ;
    if (arc_index == 1885) return "E"  ;
    if (arc_index == 1887) return "W"  ;
    if (arc_index == 1890) return "W"  ;
    if (arc_index == 1896) return "W"  ;
    if (arc_index == 1901) return "H"  ;
    if (arc_index == 1938) return "H"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 2017) return "H"  ;
    if (arc_index == 2069) return "W"  ;
    if (arc_index == 2071) return "W"  ;
    if (arc_index == 2074) return "W"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2086) return "W"  ;
    if (arc_index == 2106) return "H"  ;
    if (arc_index == 2120) return "H"  ;
    if (arc_index == 2136) return "H"  ;
    if (arc_index == 2146) return "E"  ;
    if (arc_index == 2183) return "W"  ;
    if (arc_index == 2195) return "W"  ;
    if (arc_index == 2197) return "W"  ;
    if (arc_index == 2201) return "W"  ;
    if (arc_index == 2202) return "W"  ;
    if (arc_index == 2205) return "W"  ;
    if (arc_index == 2206) return "W"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2208) return "E"  ;
    if (arc_index == 2210) return "E"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2214) return "W"  ;
    if (arc_index == 2215) return "W"  ;
    if (arc_index == 2218) return "W"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2251) return "H"  ;
    if (arc_index == 2272) return "E"  ;
    if (arc_index == 2278) return "E"  ;
    if (arc_index == 2314) return "E"  ;
    if (arc_index == 2361) return "E"  ;
    if (arc_index == 2396) return "W"  ;
    if (arc_index == 2404) return "H"  ;
    if (arc_index == 2411) return "W"  ;
    if (arc_index == 2428) return "W"  ;
    if (arc_index == 2462) return "W"  ;
    if (arc_index == 2522) return "E"  ;
    if (arc_index == 2525) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2600) return "W"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2680) return "W"  ;
    if (arc_index == 2719) return "W"  ;
    if (arc_index == 2738) return "W"  ;
    if (arc_index == 2821) return "W"  ;
    if (arc_index == 2847) return "W"  ;
    if (arc_index == 2907) return "W"  ;
    if (arc_index == 2908) return "W"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 7)) begin 
    if (arc_index == 24) return "E"  ;
    if (arc_index == 31) return "E"  ;
    if (arc_index == 91) return "E"  ;
    if (arc_index == 92) return "E"  ;
    if (arc_index == 95) return "E"  ;
    if (arc_index == 97) return "E"  ;
    if (arc_index == 101) return "E"  ;
    if (arc_index == 103) return "E"  ;
    if (arc_index == 109) return "E"  ;
    if (arc_index == 118) return "E"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 149) return "H"  ;
    if (arc_index == 156) return "H"  ;
    if (arc_index == 163) return "W"  ;
    if (arc_index == 176) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 180) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 182) return "W"  ;
    if (arc_index == 184) return "W"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 188) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 194) return "W"  ;
    if (arc_index == 229) return "W"  ;
    if (arc_index == 237) return "W"  ;
    if (arc_index == 279) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 304) return "H"  ;
    if (arc_index == 354) return "H"  ;
    if (arc_index == 359) return "H"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 420) return "E"  ;
    if (arc_index == 422) return "W"  ;
    if (arc_index == 428) return "W"  ;
    if (arc_index == 431) return "W"  ;
    if (arc_index == 433) return "W"  ;
    if (arc_index == 437) return "H"  ;
    if (arc_index == 438) return "H"  ;
    if (arc_index == 445) return "H"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 531) return "W"  ;
    if (arc_index == 532) return "H"  ;
    if (arc_index == 533) return "H"  ;
    if (arc_index == 542) return "H"  ;
    if (arc_index == 548) return "W"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 595) return "W"  ;
    if (arc_index == 616) return "W"  ;
    if (arc_index == 643) return "W"  ;
    if (arc_index == 646) return "E"  ;
    if (arc_index == 652) return "E"  ;
    if (arc_index == 658) return "H"  ;
    if (arc_index == 660) return "H"  ;
    if (arc_index == 695) return "H"  ;
    if (arc_index == 716) return "H"  ;
    if (arc_index == 729) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 742) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 759) return "W"  ;
    if (arc_index == 769) return "H"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 839) return "H"  ;
    if (arc_index == 851) return "H"  ;
    if (arc_index == 857) return "H"  ;
    if (arc_index == 898) return "E"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 969) return "E"  ;
    if (arc_index == 982) return "E"  ;
    if (arc_index == 1014) return "H"  ;
    if (arc_index == 1027) return "H"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1035) return "E"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1046) return "W"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1057) return "E"  ;
    if (arc_index == 1065) return "E"  ;
    if (arc_index == 1069) return "W"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1100) return "E"  ;
    if (arc_index == 1139) return "E"  ;
    if (arc_index == 1144) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1167) return "E"  ;
    if (arc_index == 1173) return "E"  ;
    if (arc_index == 1183) return "E"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1211) return "H"  ;
    if (arc_index == 1222) return "H"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1244) return "W"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1254) return "H"  ;
    if (arc_index == 1266) return "W"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1273) return "W"  ;
    if (arc_index == 1276) return "E"  ;
    if (arc_index == 1277) return "E"  ;
    if (arc_index == 1278) return "E"  ;
    if (arc_index == 1279) return "W"  ;
    if (arc_index == 1280) return "W"  ;
    if (arc_index == 1281) return "W"  ;
    if (arc_index == 1282) return "W"  ;
    if (arc_index == 1283) return "E"  ;
    if (arc_index == 1284) return "E"  ;
    if (arc_index == 1285) return "E"  ;
    if (arc_index == 1286) return "E"  ;
    if (arc_index == 1287) return "E"  ;
    if (arc_index == 1288) return "W"  ;
    if (arc_index == 1289) return "W"  ;
    if (arc_index == 1290) return "W"  ;
    if (arc_index == 1291) return "W"  ;
    if (arc_index == 1292) return "W"  ;
    if (arc_index == 1293) return "W"  ;
    if (arc_index == 1294) return "W"  ;
    if (arc_index == 1295) return "W"  ;
    if (arc_index == 1296) return "W"  ;
    if (arc_index == 1297) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1309) return "H"  ;
    if (arc_index == 1354) return "H"  ;
    if (arc_index == 1364) return "H"  ;
    if (arc_index == 1367) return "H"  ;
    if (arc_index == 1370) return "E"  ;
    if (arc_index == 1374) return "E"  ;
    if (arc_index == 1375) return "E"  ;
    if (arc_index == 1377) return "W"  ;
    if (arc_index == 1379) return "W"  ;
    if (arc_index == 1380) return "W"  ;
    if (arc_index == 1385) return "W"  ;
    if (arc_index == 1397) return "W"  ;
    if (arc_index == 1415) return "W"  ;
    if (arc_index == 1433) return "E"  ;
    if (arc_index == 1471) return "E"  ;
    if (arc_index == 1510) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1546) return "W"  ;
    if (arc_index == 1553) return "H"  ;
    if (arc_index == 1555) return "H"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1608) return "E"  ;
    if (arc_index == 1641) return "E"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1677) return "E"  ;
    if (arc_index == 1730) return "H"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1803) return "E"  ;
    if (arc_index == 1810) return "E"  ;
    if (arc_index == 1814) return "H"  ;
    if (arc_index == 1818) return "H"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1848) return "E"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1872) return "W"  ;
    if (arc_index == 1878) return "W"  ;
    if (arc_index == 1881) return "W"  ;
    if (arc_index == 1883) return "W"  ;
    if (arc_index == 1884) return "W"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 1900) return "E"  ;
    if (arc_index == 1923) return "H"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1976) return "W"  ;
    if (arc_index == 1988) return "W"  ;
    if (arc_index == 2010) return "W"  ;
    if (arc_index == 2019) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2039) return "H"  ;
    if (arc_index == 2042) return "H"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2077) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2087) return "W"  ;
    if (arc_index == 2128) return "H"  ;
    if (arc_index == 2130) return "E"  ;
    if (arc_index == 2133) return "E"  ;
    if (arc_index == 2141) return "E"  ;
    if (arc_index == 2142) return "H"  ;
    if (arc_index == 2147) return "E"  ;
    if (arc_index == 2201) return "E"  ;
    if (arc_index == 2206) return "E"  ;
    if (arc_index == 2220) return "E"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2251) return "E"  ;
    if (arc_index == 2263) return "E"  ;
    if (arc_index == 2270) return "E"  ;
    if (arc_index == 2273) return "H"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2316) return "W"  ;
    if (arc_index == 2318) return "W"  ;
    if (arc_index == 2321) return "W"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2330) return "W"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2372) return "W"  ;
    if (arc_index == 2418) return "W"  ;
    if (arc_index == 2426) return "H"  ;
    if (arc_index == 2428) return "H"  ;
    if (arc_index == 2435) return "H"  ;
    if (arc_index == 2444) return "E"  ;
    if (arc_index == 2446) return "E"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2507) return "E"  ;
    if (arc_index == 2517) return "E"  ;
    if (arc_index == 2524) return "E"  ;
    if (arc_index == 2528) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2599) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2725) return "E"  ;
    if (arc_index == 2736) return "E"  ;
    if (arc_index == 2764) return "E"  ;
    if (arc_index == 2837) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2922) return "W"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 9)) begin 
    if (arc_index == 139) return "W"  ;
    if (arc_index == 146) return "E"  ;
    if (arc_index == 150) return "E"  ;
    if (arc_index == 171) return "H"  ;
    if (arc_index == 289) return "H"  ;
    if (arc_index == 326) return "H"  ;
    if (arc_index == 370) return "H"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 416) return "E"  ;
    if (arc_index == 425) return "E"  ;
    if (arc_index == 427) return "E"  ;
    if (arc_index == 432) return "E"  ;
    if (arc_index == 459) return "H"  ;
    if (arc_index == 467) return "H"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 554) return "H"  ;
    if (arc_index == 620) return "H"  ;
    if (arc_index == 680) return "H"  ;
    if (arc_index == 791) return "H"  ;
    if (arc_index == 860) return "E"  ;
    if (arc_index == 861) return "H"  ;
    if (arc_index == 871) return "H"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1035) return "E"  ;
    if (arc_index == 1036) return "H"  ;
    if (arc_index == 1039) return "H"  ;
    if (arc_index == 1040) return "H"  ;
    if (arc_index == 1041) return "W"  ;
    if (arc_index == 1043) return "W"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1046) return "W"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1123) return "W"  ;
    if (arc_index == 1126) return "W"  ;
    if (arc_index == 1129) return "W"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1135) return "W"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1139) return "W"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1233) return "H"  ;
    if (arc_index == 1248) return "H"  ;
    if (arc_index == 1276) return "H"  ;
    if (arc_index == 1298) return "H"  ;
    if (arc_index == 1299) return "W"  ;
    if (arc_index == 1300) return "E"  ;
    if (arc_index == 1301) return "E"  ;
    if (arc_index == 1302) return "E"  ;
    if (arc_index == 1303) return "E"  ;
    if (arc_index == 1304) return "E"  ;
    if (arc_index == 1305) return "E"  ;
    if (arc_index == 1306) return "E"  ;
    if (arc_index == 1307) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1309) return "W"  ;
    if (arc_index == 1310) return "W"  ;
    if (arc_index == 1311) return "E"  ;
    if (arc_index == 1312) return "W"  ;
    if (arc_index == 1313) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1315) return "W"  ;
    if (arc_index == 1316) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1331) return "H"  ;
    if (arc_index == 1342) return "H"  ;
    if (arc_index == 1376) return "H"  ;
    if (arc_index == 1566) return "H"  ;
    if (arc_index == 1575) return "H"  ;
    if (arc_index == 1581) return "H"  ;
    if (arc_index == 1582) return "W"  ;
    if (arc_index == 1752) return "H"  ;
    if (arc_index == 1801) return "H"  ;
    if (arc_index == 1836) return "H"  ;
    if (arc_index == 1885) return "E"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 1900) return "E"  ;
    if (arc_index == 1945) return "H"  ;
    if (arc_index == 1974) return "E"  ;
    if (arc_index == 1988) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2061) return "H"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2119) return "E"  ;
    if (arc_index == 2150) return "H"  ;
    if (arc_index == 2164) return "H"  ;
    if (arc_index == 2178) return "W"  ;
    if (arc_index == 2180) return "W"  ;
    if (arc_index == 2203) return "E"  ;
    if (arc_index == 2211) return "E"  ;
    if (arc_index == 2272) return "E"  ;
    if (arc_index == 2295) return "H"  ;
    if (arc_index == 2325) return "H"  ;
    if (arc_index == 2377) return "W"  ;
    if (arc_index == 2448) return "H"  ;
    if (arc_index == 2455) return "H"  ;
    if (arc_index == 2575) return "H"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2654) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2726) return "W"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 9)) begin 
    if (arc_index == 8) return "W"  ;
    if (arc_index == 10) return "W"  ;
    if (arc_index == 15) return "W"  ;
    if (arc_index == 53) return "W"  ;
    if (arc_index == 56) return "W"  ;
    if (arc_index == 75) return "W"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 97) return "E"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 157) return "E"  ;
    if (arc_index == 168) return "E"  ;
    if (arc_index == 177) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 193) return "H"  ;
    if (arc_index == 196) return "H"  ;
    if (arc_index == 264) return "H"  ;
    if (arc_index == 266) return "H"  ;
    if (arc_index == 267) return "H"  ;
    if (arc_index == 272) return "H"  ;
    if (arc_index == 280) return "H"  ;
    if (arc_index == 301) return "H"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 324) return "W"  ;
    if (arc_index == 326) return "W"  ;
    if (arc_index == 332) return "E"  ;
    if (arc_index == 339) return "E"  ;
    if (arc_index == 341) return "E"  ;
    if (arc_index == 348) return "H"  ;
    if (arc_index == 425) return "H"  ;
    if (arc_index == 432) return "H"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 481) return "H"  ;
    if (arc_index == 489) return "H"  ;
    if (arc_index == 528) return "H"  ;
    if (arc_index == 529) return "E"  ;
    if (arc_index == 536) return "E"  ;
    if (arc_index == 549) return "W"  ;
    if (arc_index == 566) return "E"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 576) return "H"  ;
    if (arc_index == 590) return "H"  ;
    if (arc_index == 595) return "W"  ;
    if (arc_index == 596) return "W"  ;
    if (arc_index == 599) return "W"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 603) return "W"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 606) return "W"  ;
    if (arc_index == 607) return "W"  ;
    if (arc_index == 608) return "W"  ;
    if (arc_index == 609) return "W"  ;
    if (arc_index == 610) return "W"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 613) return "W"  ;
    if (arc_index == 622) return "W"  ;
    if (arc_index == 685) return "W"  ;
    if (arc_index == 701) return "E"  ;
    if (arc_index == 702) return "H"  ;
    if (arc_index == 704) return "H"  ;
    if (arc_index == 725) return "H"  ;
    if (arc_index == 737) return "E"  ;
    if (arc_index == 741) return "E"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 813) return "H"  ;
    if (arc_index == 817) return "H"  ;
    if (arc_index == 818) return "H"  ;
    if (arc_index == 823) return "H"  ;
    if (arc_index == 825) return "H"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 883) return "H"  ;
    if (arc_index == 975) return "H"  ;
    if (arc_index == 1034) return "W"  ;
    if (arc_index == 1037) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1058) return "H"  ;
    if (arc_index == 1066) return "H"  ;
    if (arc_index == 1067) return "E"  ;
    if (arc_index == 1071) return "E"  ;
    if (arc_index == 1133) return "W"  ;
    if (arc_index == 1142) return "W"  ;
    if (arc_index == 1205) return "W"  ;
    if (arc_index == 1251) return "W"  ;
    if (arc_index == 1253) return "W"  ;
    if (arc_index == 1255) return "H"  ;
    if (arc_index == 1268) return "H"  ;
    if (arc_index == 1298) return "H"  ;
    if (arc_index == 1316) return "H"  ;
    if (arc_index == 1320) return "E"  ;
    if (arc_index == 1321) return "W"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1323) return "W"  ;
    if (arc_index == 1324) return "W"  ;
    if (arc_index == 1325) return "W"  ;
    if (arc_index == 1326) return "E"  ;
    if (arc_index == 1327) return "W"  ;
    if (arc_index == 1328) return "W"  ;
    if (arc_index == 1329) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1331) return "W"  ;
    if (arc_index == 1332) return "W"  ;
    if (arc_index == 1333) return "W"  ;
    if (arc_index == 1334) return "W"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1338) return "W"  ;
    if (arc_index == 1339) return "E"  ;
    if (arc_index == 1340) return "E"  ;
    if (arc_index == 1341) return "W"  ;
    if (arc_index == 1353) return "H"  ;
    if (arc_index == 1354) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1363) return "W"  ;
    if (arc_index == 1375) return "W"  ;
    if (arc_index == 1382) return "W"  ;
    if (arc_index == 1394) return "W"  ;
    if (arc_index == 1398) return "H"  ;
    if (arc_index == 1399) return "H"  ;
    if (arc_index == 1426) return "H"  ;
    if (arc_index == 1460) return "E"  ;
    if (arc_index == 1475) return "E"  ;
    if (arc_index == 1479) return "E"  ;
    if (arc_index == 1544) return "W"  ;
    if (arc_index == 1554) return "W"  ;
    if (arc_index == 1577) return "W"  ;
    if (arc_index == 1583) return "W"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1597) return "H"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1654) return "E"  ;
    if (arc_index == 1682) return "E"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1769) return "E"  ;
    if (arc_index == 1770) return "E"  ;
    if (arc_index == 1774) return "H"  ;
    if (arc_index == 1780) return "H"  ;
    if (arc_index == 1797) return "H"  ;
    if (arc_index == 1806) return "E"  ;
    if (arc_index == 1858) return "H"  ;
    if (arc_index == 1869) return "E"  ;
    if (arc_index == 1880) return "E"  ;
    if (arc_index == 1907) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1967) return "H"  ;
    if (arc_index == 2068) return "H"  ;
    if (arc_index == 2070) return "H"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2081) return "W"  ;
    if (arc_index == 2083) return "H"  ;
    if (arc_index == 2100) return "H"  ;
    if (arc_index == 2141) return "H"  ;
    if (arc_index == 2172) return "H"  ;
    if (arc_index == 2186) return "H"  ;
    if (arc_index == 2267) return "H"  ;
    if (arc_index == 2286) return "H"  ;
    if (arc_index == 2295) return "H"  ;
    if (arc_index == 2303) return "E"  ;
    if (arc_index == 2310) return "E"  ;
    if (arc_index == 2317) return "H"  ;
    if (arc_index == 2320) return "W"  ;
    if (arc_index == 2326) return "W"  ;
    if (arc_index == 2329) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2333) return "W"  ;
    if (arc_index == 2343) return "W"  ;
    if (arc_index == 2345) return "E"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2351) return "W"  ;
    if (arc_index == 2358) return "W"  ;
    if (arc_index == 2361) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2386) return "W"  ;
    if (arc_index == 2389) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2403) return "W"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2407) return "W"  ;
    if (arc_index == 2410) return "W"  ;
    if (arc_index == 2413) return "W"  ;
    if (arc_index == 2415) return "W"  ;
    if (arc_index == 2419) return "W"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2470) return "H"  ;
    if (arc_index == 2476) return "H"  ;
    if (arc_index == 2482) return "H"  ;
    if (arc_index == 2537) return "E"  ;
    if (arc_index == 2548) return "E"  ;
    if (arc_index == 2599) return "W"  ;
    if (arc_index == 2606) return "W"  ;
    if (arc_index == 2615) return "W"  ;
    if (arc_index == 2643) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2689) return "E"  ;
    if (arc_index == 2690) return "E"  ;
    if (arc_index == 2696) return "E"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2775) return "W"  ;
    if (arc_index == 2776) return "E"  ;
    if (arc_index == 2825) return "E"  ;
    if (arc_index == 2830) return "E"  ;
    if (arc_index == 2831) return "E"  ;
    if (arc_index == 2836) return "E"  ;
    if (arc_index == 2895) return "E"  ;
    if (arc_index == 2902) return "E"  ;
    if (arc_index == 2904) return "W"  ;
    if (arc_index == 2907) return "W"  ;
    if (arc_index == 2913) return "W"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 10)) begin 
    if (arc_index == 11) return "E"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 197) return "E"  ;
    if (arc_index == 215) return "H"  ;
    if (arc_index == 254) return "H"  ;
    if (arc_index == 255) return "E"  ;
    if (arc_index == 267) return "E"  ;
    if (arc_index == 286) return "E"  ;
    if (arc_index == 300) return "E"  ;
    if (arc_index == 308) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 313) return "W"  ;
    if (arc_index == 316) return "W"  ;
    if (arc_index == 318) return "W"  ;
    if (arc_index == 319) return "W"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 324) return "W"  ;
    if (arc_index == 326) return "W"  ;
    if (arc_index == 327) return "W"  ;
    if (arc_index == 341) return "W"  ;
    if (arc_index == 370) return "H"  ;
    if (arc_index == 432) return "E"  ;
    if (arc_index == 503) return "H"  ;
    if (arc_index == 511) return "H"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 563) return "E"  ;
    if (arc_index == 568) return "E"  ;
    if (arc_index == 594) return "E"  ;
    if (arc_index == 598) return "H"  ;
    if (arc_index == 601) return "W"  ;
    if (arc_index == 619) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 627) return "W"  ;
    if (arc_index == 635) return "W"  ;
    if (arc_index == 639) return "W"  ;
    if (arc_index == 704) return "W"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 707) return "W"  ;
    if (arc_index == 709) return "E"  ;
    if (arc_index == 714) return "E"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 718) return "W"  ;
    if (arc_index == 723) return "W"  ;
    if (arc_index == 724) return "H"  ;
    if (arc_index == 725) return "H"  ;
    if (arc_index == 737) return "H"  ;
    if (arc_index == 824) return "H"  ;
    if (arc_index == 830) return "E"  ;
    if (arc_index == 835) return "H"  ;
    if (arc_index == 844) return "E"  ;
    if (arc_index == 905) return "H"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 1071) return "E"  ;
    if (arc_index == 1080) return "H"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1146) return "W"  ;
    if (arc_index == 1154) return "E"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1158) return "W"  ;
    if (arc_index == 1160) return "W"  ;
    if (arc_index == 1242) return "W"  ;
    if (arc_index == 1277) return "H"  ;
    if (arc_index == 1305) return "H"  ;
    if (arc_index == 1320) return "H"  ;
    if (arc_index == 1342) return "H"  ;
    if (arc_index == 1343) return "W"  ;
    if (arc_index == 1344) return "W"  ;
    if (arc_index == 1345) return "W"  ;
    if (arc_index == 1346) return "W"  ;
    if (arc_index == 1347) return "W"  ;
    if (arc_index == 1348) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1351) return "W"  ;
    if (arc_index == 1352) return "W"  ;
    if (arc_index == 1353) return "W"  ;
    if (arc_index == 1354) return "W"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1357) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1359) return "W"  ;
    if (arc_index == 1360) return "W"  ;
    if (arc_index == 1361) return "W"  ;
    if (arc_index == 1362) return "W"  ;
    if (arc_index == 1363) return "W"  ;
    if (arc_index == 1375) return "H"  ;
    if (arc_index == 1404) return "E"  ;
    if (arc_index == 1420) return "H"  ;
    if (arc_index == 1482) return "E"  ;
    if (arc_index == 1491) return "E"  ;
    if (arc_index == 1547) return "E"  ;
    if (arc_index == 1548) return "E"  ;
    if (arc_index == 1552) return "W"  ;
    if (arc_index == 1570) return "W"  ;
    if (arc_index == 1619) return "H"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1796) return "H"  ;
    if (arc_index == 1880) return "H"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1989) return "H"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2101) return "E"  ;
    if (arc_index == 2105) return "H"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2194) return "H"  ;
    if (arc_index == 2196) return "W"  ;
    if (arc_index == 2198) return "W"  ;
    if (arc_index == 2208) return "H"  ;
    if (arc_index == 2286) return "E"  ;
    if (arc_index == 2339) return "H"  ;
    if (arc_index == 2379) return "W"  ;
    if (arc_index == 2380) return "W"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2395) return "W"  ;
    if (arc_index == 2403) return "W"  ;
    if (arc_index == 2467) return "E"  ;
    if (arc_index == 2492) return "H"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2596) return "E"  ;
    if (arc_index == 2634) return "W"  ;
    if (arc_index == 2727) return "W"  ;
    if (arc_index == 2833) return "W"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2882) return "E"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2904) return "W"  ;
    if (arc_index == 2909) return "W"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2912) return "W"  ;
    if (arc_index == 2915) return "W"  ;
    if (arc_index == 2918) return "W"  ;
    if (arc_index == 2919) return "W"  ;
    if (arc_index == 2922) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 7)) begin 
    if (arc_index == 108) return "E"  ;
    if (arc_index == 139) return "E"  ;
    if (arc_index == 146) return "E"  ;
    if (arc_index == 147) return "E"  ;
    if (arc_index == 150) return "E"  ;
    if (arc_index == 237) return "H"  ;
    if (arc_index == 240) return "W"  ;
    if (arc_index == 392) return "H"  ;
    if (arc_index == 396) return "H"  ;
    if (arc_index == 421) return "W"  ;
    if (arc_index == 525) return "H"  ;
    if (arc_index == 533) return "H"  ;
    if (arc_index == 620) return "H"  ;
    if (arc_index == 661) return "E"  ;
    if (arc_index == 680) return "E"  ;
    if (arc_index == 727) return "W"  ;
    if (arc_index == 728) return "W"  ;
    if (arc_index == 732) return "W"  ;
    if (arc_index == 738) return "W"  ;
    if (arc_index == 746) return "H"  ;
    if (arc_index == 804) return "E"  ;
    if (arc_index == 857) return "H"  ;
    if (arc_index == 860) return "E"  ;
    if (arc_index == 861) return "E"  ;
    if (arc_index == 864) return "E"  ;
    if (arc_index == 867) return "E"  ;
    if (arc_index == 871) return "E"  ;
    if (arc_index == 872) return "E"  ;
    if (arc_index == 927) return "H"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 1003) return "E"  ;
    if (arc_index == 1043) return "W"  ;
    if (arc_index == 1102) return "H"  ;
    if (arc_index == 1129) return "W"  ;
    if (arc_index == 1135) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1180) return "E"  ;
    if (arc_index == 1248) return "W"  ;
    if (arc_index == 1258) return "W"  ;
    if (arc_index == 1299) return "H"  ;
    if (arc_index == 1307) return "W"  ;
    if (arc_index == 1342) return "H"  ;
    if (arc_index == 1364) return "H"  ;
    if (arc_index == 1365) return "H"  ;
    if (arc_index == 1366) return "H"  ;
    if (arc_index == 1367) return "H"  ;
    if (arc_index == 1368) return "H"  ;
    if (arc_index == 1369) return "E"  ;
    if (arc_index == 1370) return "E"  ;
    if (arc_index == 1371) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1373) return "E"  ;
    if (arc_index == 1374) return "E"  ;
    if (arc_index == 1375) return "E"  ;
    if (arc_index == 1376) return "E"  ;
    if (arc_index == 1377) return "E"  ;
    if (arc_index == 1378) return "W"  ;
    if (arc_index == 1379) return "W"  ;
    if (arc_index == 1380) return "W"  ;
    if (arc_index == 1381) return "W"  ;
    if (arc_index == 1382) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1384) return "W"  ;
    if (arc_index == 1385) return "W"  ;
    if (arc_index == 1397) return "H"  ;
    if (arc_index == 1442) return "H"  ;
    if (arc_index == 1513) return "E"  ;
    if (arc_index == 1563) return "E"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1565) return "W"  ;
    if (arc_index == 1568) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1641) return "H"  ;
    if (arc_index == 1723) return "E"  ;
    if (arc_index == 1818) return "H"  ;
    if (arc_index == 1902) return "H"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2011) return "H"  ;
    if (arc_index == 2016) return "E"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2086) return "W"  ;
    if (arc_index == 2127) return "H"  ;
    if (arc_index == 2195) return "W"  ;
    if (arc_index == 2216) return "H"  ;
    if (arc_index == 2230) return "H"  ;
    if (arc_index == 2314) return "W"  ;
    if (arc_index == 2361) return "H"  ;
    if (arc_index == 2514) return "H"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2657) return "W"  ;
    if (arc_index == 2660) return "W"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2813) return "E"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 5)) begin 
    if (arc_index == 4) return "W"  ;
    if (arc_index == 86) return "E"  ;
    if (arc_index == 95) return "W"  ;
    if (arc_index == 164) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 247) return "W"  ;
    if (arc_index == 248) return "W"  ;
    if (arc_index == 251) return "W"  ;
    if (arc_index == 256) return "W"  ;
    if (arc_index == 259) return "H"  ;
    if (arc_index == 262) return "W"  ;
    if (arc_index == 263) return "W"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 311) return "W"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 340) return "W"  ;
    if (arc_index == 414) return "H"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 547) return "H"  ;
    if (arc_index == 550) return "H"  ;
    if (arc_index == 555) return "H"  ;
    if (arc_index == 571) return "H"  ;
    if (arc_index == 577) return "H"  ;
    if (arc_index == 642) return "H"  ;
    if (arc_index == 683) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 749) return "E"  ;
    if (arc_index == 760) return "E"  ;
    if (arc_index == 762) return "E"  ;
    if (arc_index == 763) return "E"  ;
    if (arc_index == 765) return "E"  ;
    if (arc_index == 768) return "H"  ;
    if (arc_index == 772) return "H"  ;
    if (arc_index == 780) return "E"  ;
    if (arc_index == 782) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 826) return "W"  ;
    if (arc_index == 843) return "W"  ;
    if (arc_index == 879) return "H"  ;
    if (arc_index == 889) return "E"  ;
    if (arc_index == 949) return "H"  ;
    if (arc_index == 1076) return "H"  ;
    if (arc_index == 1120) return "W"  ;
    if (arc_index == 1124) return "H"  ;
    if (arc_index == 1187) return "H"  ;
    if (arc_index == 1257) return "H"  ;
    if (arc_index == 1286) return "W"  ;
    if (arc_index == 1321) return "H"  ;
    if (arc_index == 1364) return "H"  ;
    if (arc_index == 1386) return "H"  ;
    if (arc_index == 1387) return "E"  ;
    if (arc_index == 1388) return "W"  ;
    if (arc_index == 1389) return "W"  ;
    if (arc_index == 1390) return "W"  ;
    if (arc_index == 1391) return "W"  ;
    if (arc_index == 1392) return "E"  ;
    if (arc_index == 1393) return "E"  ;
    if (arc_index == 1394) return "E"  ;
    if (arc_index == 1395) return "W"  ;
    if (arc_index == 1396) return "W"  ;
    if (arc_index == 1397) return "W"  ;
    if (arc_index == 1398) return "W"  ;
    if (arc_index == 1399) return "W"  ;
    if (arc_index == 1400) return "W"  ;
    if (arc_index == 1401) return "W"  ;
    if (arc_index == 1402) return "E"  ;
    if (arc_index == 1403) return "E"  ;
    if (arc_index == 1404) return "E"  ;
    if (arc_index == 1405) return "E"  ;
    if (arc_index == 1406) return "W"  ;
    if (arc_index == 1407) return "W"  ;
    if (arc_index == 1408) return "W"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1419) return "H"  ;
    if (arc_index == 1432) return "H"  ;
    if (arc_index == 1441) return "H"  ;
    if (arc_index == 1453) return "H"  ;
    if (arc_index == 1454) return "W"  ;
    if (arc_index == 1459) return "W"  ;
    if (arc_index == 1463) return "W"  ;
    if (arc_index == 1464) return "H"  ;
    if (arc_index == 1465) return "H"  ;
    if (arc_index == 1466) return "H"  ;
    if (arc_index == 1473) return "H"  ;
    if (arc_index == 1580) return "H"  ;
    if (arc_index == 1663) return "H"  ;
    if (arc_index == 1672) return "H"  ;
    if (arc_index == 1694) return "H"  ;
    if (arc_index == 1696) return "H"  ;
    if (arc_index == 1697) return "H"  ;
    if (arc_index == 1698) return "H"  ;
    if (arc_index == 1699) return "H"  ;
    if (arc_index == 1702) return "H"  ;
    if (arc_index == 1703) return "H"  ;
    if (arc_index == 1707) return "H"  ;
    if (arc_index == 1710) return "H"  ;
    if (arc_index == 1738) return "E"  ;
    if (arc_index == 1757) return "E"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1761) return "E"  ;
    if (arc_index == 1800) return "W"  ;
    if (arc_index == 1816) return "W"  ;
    if (arc_index == 1838) return "W"  ;
    if (arc_index == 1840) return "H"  ;
    if (arc_index == 1854) return "E"  ;
    if (arc_index == 1866) return "W"  ;
    if (arc_index == 1924) return "H"  ;
    if (arc_index == 1990) return "E"  ;
    if (arc_index == 2025) return "E"  ;
    if (arc_index == 2026) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2033) return "H"  ;
    if (arc_index == 2041) return "E"  ;
    if (arc_index == 2096) return "E"  ;
    if (arc_index == 2149) return "H"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2223) return "E"  ;
    if (arc_index == 2238) return "H"  ;
    if (arc_index == 2252) return "H"  ;
    if (arc_index == 2265) return "H"  ;
    if (arc_index == 2290) return "W"  ;
    if (arc_index == 2291) return "W"  ;
    if (arc_index == 2297) return "W"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2301) return "W"  ;
    if (arc_index == 2305) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2383) return "H"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2487) return "W"  ;
    if (arc_index == 2501) return "W"  ;
    if (arc_index == 2530) return "W"  ;
    if (arc_index == 2536) return "H"  ;
    if (arc_index == 2544) return "H"  ;
    if (arc_index == 2546) return "H"  ;
    if (arc_index == 2559) return "H"  ;
    if (arc_index == 2563) return "H"  ;
    if (arc_index == 2565) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2604) return "W"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2731) return "E"  ;
    if (arc_index == 2732) return "E"  ;
    if (arc_index == 2742) return "E"  ;
    if (arc_index == 2744) return "E"  ;
    if (arc_index == 2749) return "E"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2779) return "E"  ;
    if (arc_index == 2782) return "E"  ;
    if (arc_index == 2786) return "E"  ;
    if (arc_index == 2790) return "E"  ;
    if (arc_index == 2816) return "W"  ;
    if (arc_index == 2829) return "W"  ;
    if (arc_index == 2835) return "W"  ;
    if (arc_index == 2839) return "W"  ;
    if (arc_index == 2841) return "W"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2849) return "E"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2864) return "E"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2873) return "E"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 6)) begin 
    if (arc_index == 113) return "E"  ;
    if (arc_index == 281) return "H"  ;
    if (arc_index == 436) return "H"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 550) return "W"  ;
    if (arc_index == 553) return "W"  ;
    if (arc_index == 555) return "W"  ;
    if (arc_index == 559) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 565) return "W"  ;
    if (arc_index == 567) return "W"  ;
    if (arc_index == 569) return "H"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 571) return "W"  ;
    if (arc_index == 577) return "H"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 664) return "H"  ;
    if (arc_index == 698) return "W"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 712) return "W"  ;
    if (arc_index == 722) return "W"  ;
    if (arc_index == 788) return "E"  ;
    if (arc_index == 790) return "H"  ;
    if (arc_index == 855) return "W"  ;
    if (arc_index == 863) return "W"  ;
    if (arc_index == 901) return "H"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 971) return "H"  ;
    if (arc_index == 1146) return "H"  ;
    if (arc_index == 1197) return "E"  ;
    if (arc_index == 1343) return "H"  ;
    if (arc_index == 1386) return "H"  ;
    if (arc_index == 1408) return "W"  ;
    if (arc_index == 1409) return "E"  ;
    if (arc_index == 1410) return "E"  ;
    if (arc_index == 1411) return "E"  ;
    if (arc_index == 1412) return "E"  ;
    if (arc_index == 1413) return "E"  ;
    if (arc_index == 1414) return "E"  ;
    if (arc_index == 1415) return "E"  ;
    if (arc_index == 1416) return "E"  ;
    if (arc_index == 1417) return "W"  ;
    if (arc_index == 1418) return "W"  ;
    if (arc_index == 1419) return "W"  ;
    if (arc_index == 1420) return "E"  ;
    if (arc_index == 1421) return "E"  ;
    if (arc_index == 1422) return "E"  ;
    if (arc_index == 1423) return "E"  ;
    if (arc_index == 1424) return "W"  ;
    if (arc_index == 1425) return "W"  ;
    if (arc_index == 1426) return "E"  ;
    if (arc_index == 1427) return "E"  ;
    if (arc_index == 1428) return "E"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1441) return "H"  ;
    if (arc_index == 1472) return "E"  ;
    if (arc_index == 1486) return "H"  ;
    if (arc_index == 1498) return "E"  ;
    if (arc_index == 1685) return "H"  ;
    if (arc_index == 1695) return "E"  ;
    if (arc_index == 1700) return "E"  ;
    if (arc_index == 1701) return "E"  ;
    if (arc_index == 1704) return "E"  ;
    if (arc_index == 1705) return "E"  ;
    if (arc_index == 1708) return "E"  ;
    if (arc_index == 1714) return "E"  ;
    if (arc_index == 1761) return "W"  ;
    if (arc_index == 1762) return "W"  ;
    if (arc_index == 1767) return "W"  ;
    if (arc_index == 1771) return "W"  ;
    if (arc_index == 1772) return "W"  ;
    if (arc_index == 1838) return "E"  ;
    if (arc_index == 1862) return "H"  ;
    if (arc_index == 1946) return "H"  ;
    if (arc_index == 1971) return "W"  ;
    if (arc_index == 2025) return "E"  ;
    if (arc_index == 2037) return "E"  ;
    if (arc_index == 2055) return "H"  ;
    if (arc_index == 2094) return "W"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2102) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2110) return "W"  ;
    if (arc_index == 2171) return "H"  ;
    if (arc_index == 2260) return "H"  ;
    if (arc_index == 2274) return "H"  ;
    if (arc_index == 2335) return "W"  ;
    if (arc_index == 2341) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2405) return "H"  ;
    if (arc_index == 2544) return "E"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2558) return "H"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2732) return "E"  ;
    if (arc_index == 2737) return "E"  ;
    if (arc_index == 2776) return "E"  ;
    if (arc_index == 2777) return "E"  ;
    if (arc_index == 2791) return "E"  ;
    if (arc_index == 2853) return "E"  ;
    if (arc_index == 2858) return "E"  ;
    if (arc_index == 2916) return "W"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 5)) begin 
    if (arc_index == 0) return "W"  ;
    if (arc_index == 1) return "W"  ;
    if (arc_index == 3) return "W"  ;
    if (arc_index == 30) return "W"  ;
    if (arc_index == 33) return "E"  ;
    if (arc_index == 38) return "E"  ;
    if (arc_index == 43) return "E"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 52) return "E"  ;
    if (arc_index == 53) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 57) return "E"  ;
    if (arc_index == 62) return "E"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 68) return "E"  ;
    if (arc_index == 72) return "E"  ;
    if (arc_index == 106) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 116) return "W"  ;
    if (arc_index == 123) return "W"  ;
    if (arc_index == 125) return "W"  ;
    if (arc_index == 128) return "E"  ;
    if (arc_index == 130) return "E"  ;
    if (arc_index == 159) return "W"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 210) return "W"  ;
    if (arc_index == 222) return "W"  ;
    if (arc_index == 227) return "W"  ;
    if (arc_index == 238) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 303) return "H"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 336) return "W"  ;
    if (arc_index == 343) return "W"  ;
    if (arc_index == 346) return "W"  ;
    if (arc_index == 349) return "W"  ;
    if (arc_index == 350) return "W"  ;
    if (arc_index == 362) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 367) return "W"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 399) return "E"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 412) return "W"  ;
    if (arc_index == 414) return "W"  ;
    if (arc_index == 447) return "W"  ;
    if (arc_index == 458) return "H"  ;
    if (arc_index == 467) return "H"  ;
    if (arc_index == 474) return "H"  ;
    if (arc_index == 490) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 497) return "E"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 530) return "W"  ;
    if (arc_index == 540) return "W"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 591) return "H"  ;
    if (arc_index == 599) return "H"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 663) return "W"  ;
    if (arc_index == 674) return "E"  ;
    if (arc_index == 686) return "H"  ;
    if (arc_index == 691) return "W"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 726) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 757) return "W"  ;
    if (arc_index == 759) return "W"  ;
    if (arc_index == 769) return "E"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 812) return "H"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 862) return "W"  ;
    if (arc_index == 879) return "W"  ;
    if (arc_index == 904) return "E"  ;
    if (arc_index == 923) return "H"  ;
    if (arc_index == 928) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 971) return "E"  ;
    if (arc_index == 972) return "W"  ;
    if (arc_index == 973) return "E"  ;
    if (arc_index == 974) return "E"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 980) return "E"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 983) return "E"  ;
    if (arc_index == 985) return "E"  ;
    if (arc_index == 986) return "E"  ;
    if (arc_index == 987) return "W"  ;
    if (arc_index == 988) return "W"  ;
    if (arc_index == 991) return "W"  ;
    if (arc_index == 993) return "H"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1096) return "W"  ;
    if (arc_index == 1168) return "H"  ;
    if (arc_index == 1195) return "H"  ;
    if (arc_index == 1196) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1214) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1269) return "E"  ;
    if (arc_index == 1279) return "E"  ;
    if (arc_index == 1281) return "E"  ;
    if (arc_index == 1292) return "W"  ;
    if (arc_index == 1296) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1325) return "W"  ;
    if (arc_index == 1365) return "H"  ;
    if (arc_index == 1368) return "H"  ;
    if (arc_index == 1385) return "H"  ;
    if (arc_index == 1393) return "H"  ;
    if (arc_index == 1408) return "H"  ;
    if (arc_index == 1422) return "H"  ;
    if (arc_index == 1430) return "H"  ;
    if (arc_index == 1431) return "H"  ;
    if (arc_index == 1432) return "H"  ;
    if (arc_index == 1433) return "H"  ;
    if (arc_index == 1434) return "E"  ;
    if (arc_index == 1435) return "E"  ;
    if (arc_index == 1436) return "E"  ;
    if (arc_index == 1437) return "W"  ;
    if (arc_index == 1438) return "W"  ;
    if (arc_index == 1439) return "W"  ;
    if (arc_index == 1440) return "W"  ;
    if (arc_index == 1441) return "W"  ;
    if (arc_index == 1442) return "W"  ;
    if (arc_index == 1443) return "E"  ;
    if (arc_index == 1444) return "W"  ;
    if (arc_index == 1445) return "E"  ;
    if (arc_index == 1446) return "E"  ;
    if (arc_index == 1447) return "E"  ;
    if (arc_index == 1448) return "W"  ;
    if (arc_index == 1449) return "E"  ;
    if (arc_index == 1450) return "E"  ;
    if (arc_index == 1451) return "E"  ;
    if (arc_index == 1462) return "W"  ;
    if (arc_index == 1463) return "H"  ;
    if (arc_index == 1470) return "H"  ;
    if (arc_index == 1498) return "H"  ;
    if (arc_index == 1508) return "H"  ;
    if (arc_index == 1514) return "H"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1522) return "E"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1615) return "W"  ;
    if (arc_index == 1621) return "W"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1635) return "E"  ;
    if (arc_index == 1648) return "E"  ;
    if (arc_index == 1707) return "H"  ;
    if (arc_index == 1710) return "H"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1773) return "E"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1802) return "W"  ;
    if (arc_index == 1821) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1855) return "W"  ;
    if (arc_index == 1864) return "W"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1881) return "W"  ;
    if (arc_index == 1883) return "W"  ;
    if (arc_index == 1884) return "H"  ;
    if (arc_index == 1900) return "E"  ;
    if (arc_index == 1902) return "E"  ;
    if (arc_index == 1909) return "E"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1968) return "H"  ;
    if (arc_index == 1973) return "H"  ;
    if (arc_index == 2004) return "E"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2048) return "E"  ;
    if (arc_index == 2061) return "E"  ;
    if (arc_index == 2077) return "H"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2112) return "W"  ;
    if (arc_index == 2113) return "E"  ;
    if (arc_index == 2117) return "E"  ;
    if (arc_index == 2118) return "E"  ;
    if (arc_index == 2119) return "E"  ;
    if (arc_index == 2120) return "E"  ;
    if (arc_index == 2127) return "E"  ;
    if (arc_index == 2128) return "E"  ;
    if (arc_index == 2130) return "E"  ;
    if (arc_index == 2133) return "E"  ;
    if (arc_index == 2145) return "E"  ;
    if (arc_index == 2156) return "E"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2169) return "E"  ;
    if (arc_index == 2174) return "E"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2189) return "W"  ;
    if (arc_index == 2190) return "W"  ;
    if (arc_index == 2193) return "H"  ;
    if (arc_index == 2202) return "H"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2259) return "W"  ;
    if (arc_index == 2275) return "W"  ;
    if (arc_index == 2279) return "W"  ;
    if (arc_index == 2281) return "W"  ;
    if (arc_index == 2282) return "H"  ;
    if (arc_index == 2283) return "W"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2296) return "H"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2425) return "E"  ;
    if (arc_index == 2427) return "H"  ;
    if (arc_index == 2430) return "H"  ;
    if (arc_index == 2449) return "H"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2491) return "E"  ;
    if (arc_index == 2493) return "E"  ;
    if (arc_index == 2498) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2533) return "W"  ;
    if (arc_index == 2534) return "E"  ;
    if (arc_index == 2551) return "W"  ;
    if (arc_index == 2580) return "H"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2708) return "W"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2752) return "E"  ;
    if (arc_index == 2764) return "E"  ;
    if (arc_index == 2767) return "E"  ;
    if (arc_index == 2771) return "E"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2841) return "E"  ;
    if (arc_index == 2905) return "W"  ;
    if (arc_index == 2919) return "W"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 6)) begin 
    if (arc_index == 86) return "E"  ;
    if (arc_index == 95) return "W"  ;
    if (arc_index == 113) return "W"  ;
    if (arc_index == 164) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 247) return "W"  ;
    if (arc_index == 248) return "W"  ;
    if (arc_index == 251) return "W"  ;
    if (arc_index == 256) return "W"  ;
    if (arc_index == 259) return "W"  ;
    if (arc_index == 262) return "W"  ;
    if (arc_index == 263) return "W"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 325) return "H"  ;
    if (arc_index == 340) return "W"  ;
    if (arc_index == 436) return "W"  ;
    if (arc_index == 480) return "H"  ;
    if (arc_index == 485) return "H"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 553) return "E"  ;
    if (arc_index == 562) return "E"  ;
    if (arc_index == 613) return "H"  ;
    if (arc_index == 621) return "H"  ;
    if (arc_index == 642) return "W"  ;
    if (arc_index == 683) return "W"  ;
    if (arc_index == 698) return "W"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 708) return "H"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 722) return "W"  ;
    if (arc_index == 749) return "E"  ;
    if (arc_index == 780) return "E"  ;
    if (arc_index == 782) return "E"  ;
    if (arc_index == 834) return "H"  ;
    if (arc_index == 843) return "W"  ;
    if (arc_index == 855) return "W"  ;
    if (arc_index == 863) return "W"  ;
    if (arc_index == 889) return "E"  ;
    if (arc_index == 901) return "E"  ;
    if (arc_index == 945) return "H"  ;
    if (arc_index == 971) return "H"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1015) return "H"  ;
    if (arc_index == 1094) return "E"  ;
    if (arc_index == 1120) return "W"  ;
    if (arc_index == 1146) return "W"  ;
    if (arc_index == 1190) return "H"  ;
    if (arc_index == 1286) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1387) return "H"  ;
    if (arc_index == 1392) return "E"  ;
    if (arc_index == 1394) return "E"  ;
    if (arc_index == 1402) return "E"  ;
    if (arc_index == 1410) return "E"  ;
    if (arc_index == 1411) return "E"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1413) return "W"  ;
    if (arc_index == 1414) return "W"  ;
    if (arc_index == 1415) return "W"  ;
    if (arc_index == 1421) return "W"  ;
    if (arc_index == 1422) return "W"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1427) return "W"  ;
    if (arc_index == 1428) return "W"  ;
    if (arc_index == 1430) return "H"  ;
    if (arc_index == 1452) return "H"  ;
    if (arc_index == 1453) return "W"  ;
    if (arc_index == 1454) return "W"  ;
    if (arc_index == 1455) return "W"  ;
    if (arc_index == 1456) return "W"  ;
    if (arc_index == 1457) return "E"  ;
    if (arc_index == 1458) return "E"  ;
    if (arc_index == 1459) return "W"  ;
    if (arc_index == 1460) return "W"  ;
    if (arc_index == 1461) return "W"  ;
    if (arc_index == 1462) return "W"  ;
    if (arc_index == 1463) return "W"  ;
    if (arc_index == 1464) return "W"  ;
    if (arc_index == 1465) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1467) return "E"  ;
    if (arc_index == 1468) return "E"  ;
    if (arc_index == 1469) return "E"  ;
    if (arc_index == 1470) return "E"  ;
    if (arc_index == 1471) return "E"  ;
    if (arc_index == 1472) return "E"  ;
    if (arc_index == 1473) return "W"  ;
    if (arc_index == 1485) return "H"  ;
    if (arc_index == 1486) return "H"  ;
    if (arc_index == 1498) return "H"  ;
    if (arc_index == 1530) return "H"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1685) return "W"  ;
    if (arc_index == 1704) return "W"  ;
    if (arc_index == 1705) return "E"  ;
    if (arc_index == 1729) return "H"  ;
    if (arc_index == 1738) return "E"  ;
    if (arc_index == 1757) return "E"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1760) return "E"  ;
    if (arc_index == 1773) return "E"  ;
    if (arc_index == 1800) return "W"  ;
    if (arc_index == 1816) return "W"  ;
    if (arc_index == 1854) return "E"  ;
    if (arc_index == 1862) return "E"  ;
    if (arc_index == 1906) return "H"  ;
    if (arc_index == 1971) return "H"  ;
    if (arc_index == 1990) return "H"  ;
    if (arc_index == 2025) return "H"  ;
    if (arc_index == 2026) return "E"  ;
    if (arc_index == 2041) return "E"  ;
    if (arc_index == 2055) return "E"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2099) return "H"  ;
    if (arc_index == 2109) return "H"  ;
    if (arc_index == 2171) return "H"  ;
    if (arc_index == 2215) return "H"  ;
    if (arc_index == 2223) return "E"  ;
    if (arc_index == 2252) return "W"  ;
    if (arc_index == 2260) return "W"  ;
    if (arc_index == 2274) return "W"  ;
    if (arc_index == 2290) return "W"  ;
    if (arc_index == 2291) return "W"  ;
    if (arc_index == 2297) return "W"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2301) return "W"  ;
    if (arc_index == 2304) return "H"  ;
    if (arc_index == 2305) return "W"  ;
    if (arc_index == 2318) return "H"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2449) return "H"  ;
    if (arc_index == 2531) return "E"  ;
    if (arc_index == 2550) return "E"  ;
    if (arc_index == 2565) return "E"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2602) return "H"  ;
    if (arc_index == 2604) return "W"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2731) return "E"  ;
    if (arc_index == 2742) return "E"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2776) return "E"  ;
    if (arc_index == 2782) return "E"  ;
    if (arc_index == 2791) return "E"  ;
    if (arc_index == 2816) return "W"  ;
    if (arc_index == 2829) return "W"  ;
    if (arc_index == 2848) return "W"  ;
    if (arc_index == 2852) return "W"  ;
    if (arc_index == 2864) return "E"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2873) return "E"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 8)) begin 
    if (arc_index == 11) return "E"  ;
    if (arc_index == 30) return "E"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 161) return "E"  ;
    if (arc_index == 164) return "E"  ;
    if (arc_index == 167) return "W"  ;
    if (arc_index == 175) return "W"  ;
    if (arc_index == 177) return "W"  ;
    if (arc_index == 199) return "W"  ;
    if (arc_index == 213) return "W"  ;
    if (arc_index == 215) return "E"  ;
    if (arc_index == 220) return "E"  ;
    if (arc_index == 228) return "E"  ;
    if (arc_index == 231) return "E"  ;
    if (arc_index == 242) return "E"  ;
    if (arc_index == 249) return "E"  ;
    if (arc_index == 250) return "E"  ;
    if (arc_index == 252) return "E"  ;
    if (arc_index == 253) return "E"  ;
    if (arc_index == 255) return "E"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 260) return "W"  ;
    if (arc_index == 275) return "W"  ;
    if (arc_index == 301) return "W"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 315) return "W"  ;
    if (arc_index == 347) return "H"  ;
    if (arc_index == 354) return "H"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 420) return "E"  ;
    if (arc_index == 433) return "E"  ;
    if (arc_index == 502) return "H"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 528) return "E"  ;
    if (arc_index == 547) return "W"  ;
    if (arc_index == 566) return "E"  ;
    if (arc_index == 568) return "E"  ;
    if (arc_index == 601) return "W"  ;
    if (arc_index == 613) return "W"  ;
    if (arc_index == 619) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 635) return "H"  ;
    if (arc_index == 643) return "H"  ;
    if (arc_index == 649) return "H"  ;
    if (arc_index == 660) return "H"  ;
    if (arc_index == 685) return "E"  ;
    if (arc_index == 689) return "E"  ;
    if (arc_index == 692) return "E"  ;
    if (arc_index == 695) return "E"  ;
    if (arc_index == 700) return "E"  ;
    if (arc_index == 701) return "E"  ;
    if (arc_index == 702) return "E"  ;
    if (arc_index == 703) return "E"  ;
    if (arc_index == 713) return "E"  ;
    if (arc_index == 721) return "E"  ;
    if (arc_index == 730) return "H"  ;
    if (arc_index == 749) return "E"  ;
    if (arc_index == 814) return "E"  ;
    if (arc_index == 815) return "W"  ;
    if (arc_index == 816) return "W"  ;
    if (arc_index == 819) return "W"  ;
    if (arc_index == 821) return "W"  ;
    if (arc_index == 822) return "W"  ;
    if (arc_index == 826) return "W"  ;
    if (arc_index == 827) return "W"  ;
    if (arc_index == 831) return "W"  ;
    if (arc_index == 832) return "W"  ;
    if (arc_index == 833) return "W"  ;
    if (arc_index == 844) return "E"  ;
    if (arc_index == 856) return "H"  ;
    if (arc_index == 892) return "E"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 967) return "H"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 1037) return "H"  ;
    if (arc_index == 1040) return "W"  ;
    if (arc_index == 1070) return "E"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1091) return "E"  ;
    if (arc_index == 1118) return "E"  ;
    if (arc_index == 1136) return "E"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1212) return "H"  ;
    if (arc_index == 1236) return "W"  ;
    if (arc_index == 1239) return "W"  ;
    if (arc_index == 1251) return "W"  ;
    if (arc_index == 1259) return "W"  ;
    if (arc_index == 1263) return "W"  ;
    if (arc_index == 1316) return "W"  ;
    if (arc_index == 1329) return "W"  ;
    if (arc_index == 1344) return "W"  ;
    if (arc_index == 1345) return "W"  ;
    if (arc_index == 1348) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1359) return "W"  ;
    if (arc_index == 1362) return "W"  ;
    if (arc_index == 1404) return "E"  ;
    if (arc_index == 1409) return "H"  ;
    if (arc_index == 1410) return "H"  ;
    if (arc_index == 1414) return "H"  ;
    if (arc_index == 1421) return "E"  ;
    if (arc_index == 1426) return "E"  ;
    if (arc_index == 1445) return "E"  ;
    if (arc_index == 1452) return "H"  ;
    if (arc_index == 1461) return "E"  ;
    if (arc_index == 1474) return "E"  ;
    if (arc_index == 1475) return "E"  ;
    if (arc_index == 1476) return "W"  ;
    if (arc_index == 1477) return "W"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1479) return "W"  ;
    if (arc_index == 1480) return "W"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1482) return "E"  ;
    if (arc_index == 1483) return "W"  ;
    if (arc_index == 1484) return "W"  ;
    if (arc_index == 1485) return "W"  ;
    if (arc_index == 1486) return "W"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1488) return "W"  ;
    if (arc_index == 1489) return "W"  ;
    if (arc_index == 1490) return "W"  ;
    if (arc_index == 1491) return "E"  ;
    if (arc_index == 1492) return "W"  ;
    if (arc_index == 1493) return "E"  ;
    if (arc_index == 1494) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1501) return "W"  ;
    if (arc_index == 1507) return "H"  ;
    if (arc_index == 1544) return "W"  ;
    if (arc_index == 1552) return "H"  ;
    if (arc_index == 1583) return "H"  ;
    if (arc_index == 1613) return "E"  ;
    if (arc_index == 1619) return "E"  ;
    if (arc_index == 1653) return "E"  ;
    if (arc_index == 1666) return "E"  ;
    if (arc_index == 1679) return "E"  ;
    if (arc_index == 1685) return "E"  ;
    if (arc_index == 1688) return "E"  ;
    if (arc_index == 1705) return "E"  ;
    if (arc_index == 1708) return "E"  ;
    if (arc_index == 1751) return "H"  ;
    if (arc_index == 1763) return "H"  ;
    if (arc_index == 1775) return "H"  ;
    if (arc_index == 1778) return "W"  ;
    if (arc_index == 1791) return "W"  ;
    if (arc_index == 1796) return "E"  ;
    if (arc_index == 1797) return "E"  ;
    if (arc_index == 1811) return "E"  ;
    if (arc_index == 1825) return "E"  ;
    if (arc_index == 1852) return "E"  ;
    if (arc_index == 1928) return "H"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1964) return "E"  ;
    if (arc_index == 1978) return "E"  ;
    if (arc_index == 1989) return "E"  ;
    if (arc_index == 1996) return "E"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2012) return "H"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2072) return "W"  ;
    if (arc_index == 2090) return "W"  ;
    if (arc_index == 2091) return "W"  ;
    if (arc_index == 2098) return "W"  ;
    if (arc_index == 2100) return "E"  ;
    if (arc_index == 2106) return "E"  ;
    if (arc_index == 2108) return "E"  ;
    if (arc_index == 2121) return "H"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2198) return "W"  ;
    if (arc_index == 2214) return "W"  ;
    if (arc_index == 2237) return "H"  ;
    if (arc_index == 2295) return "E"  ;
    if (arc_index == 2326) return "H"  ;
    if (arc_index == 2329) return "H"  ;
    if (arc_index == 2340) return "H"  ;
    if (arc_index == 2342) return "W"  ;
    if (arc_index == 2344) return "W"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2364) return "W"  ;
    if (arc_index == 2367) return "W"  ;
    if (arc_index == 2379) return "W"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2424) return "W"  ;
    if (arc_index == 2471) return "H"  ;
    if (arc_index == 2484) return "H"  ;
    if (arc_index == 2490) return "H"  ;
    if (arc_index == 2492) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2600) return "E"  ;
    if (arc_index == 2601) return "E"  ;
    if (arc_index == 2611) return "W"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2624) return "H"  ;
    if (arc_index == 2634) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2753) return "E"  ;
    if (arc_index == 2768) return "E"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2776) return "E"  ;
    if (arc_index == 2818) return "E"  ;
    if (arc_index == 2830) return "E"  ;
    if (arc_index == 2833) return "E"  ;
    if (arc_index == 2836) return "E"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2882) return "E"  ;
    if (arc_index == 2901) return "E"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2915) return "W"  ;
    if (arc_index == 2918) return "W"  ;
    if (arc_index == 2919) return "W"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 5)) begin 
    if (arc_index == 27) return "W"  ;
    if (arc_index == 114) return "E"  ;
    if (arc_index == 137) return "E"  ;
    if (arc_index == 140) return "E"  ;
    if (arc_index == 143) return "E"  ;
    if (arc_index == 223) return "E"  ;
    if (arc_index == 331) return "E"  ;
    if (arc_index == 352) return "W"  ;
    if (arc_index == 355) return "W"  ;
    if (arc_index == 357) return "W"  ;
    if (arc_index == 360) return "W"  ;
    if (arc_index == 368) return "W"  ;
    if (arc_index == 369) return "H"  ;
    if (arc_index == 372) return "W"  ;
    if (arc_index == 374) return "W"  ;
    if (arc_index == 392) return "E"  ;
    if (arc_index == 397) return "E"  ;
    if (arc_index == 399) return "E"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 401) return "E"  ;
    if (arc_index == 402) return "E"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 404) return "E"  ;
    if (arc_index == 405) return "E"  ;
    if (arc_index == 406) return "E"  ;
    if (arc_index == 408) return "E"  ;
    if (arc_index == 410) return "E"  ;
    if (arc_index == 412) return "E"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 414) return "E"  ;
    if (arc_index == 415) return "E"  ;
    if (arc_index == 418) return "W"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 434) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 474) return "W"  ;
    if (arc_index == 524) return "H"  ;
    if (arc_index == 638) return "W"  ;
    if (arc_index == 657) return "H"  ;
    if (arc_index == 660) return "E"  ;
    if (arc_index == 665) return "H"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 677) return "E"  ;
    if (arc_index == 728) return "W"  ;
    if (arc_index == 752) return "H"  ;
    if (arc_index == 793) return "H"  ;
    if (arc_index == 796) return "H"  ;
    if (arc_index == 806) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 825) return "W"  ;
    if (arc_index == 850) return "W"  ;
    if (arc_index == 862) return "W"  ;
    if (arc_index == 873) return "W"  ;
    if (arc_index == 874) return "W"  ;
    if (arc_index == 878) return "H"  ;
    if (arc_index == 879) return "H"  ;
    if (arc_index == 927) return "E"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 968) return "W"  ;
    if (arc_index == 984) return "W"  ;
    if (arc_index == 989) return "H"  ;
    if (arc_index == 991) return "H"  ;
    if (arc_index == 992) return "E"  ;
    if (arc_index == 999) return "E"  ;
    if (arc_index == 1003) return "E"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1041) return "E"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1059) return "H"  ;
    if (arc_index == 1069) return "W"  ;
    if (arc_index == 1123) return "W"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1171) return "W"  ;
    if (arc_index == 1204) return "E"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1234) return "H"  ;
    if (arc_index == 1246) return "W"  ;
    if (arc_index == 1262) return "W"  ;
    if (arc_index == 1315) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1371) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1381) return "W"  ;
    if (arc_index == 1393) return "W"  ;
    if (arc_index == 1431) return "H"  ;
    if (arc_index == 1447) return "W"  ;
    if (arc_index == 1474) return "H"  ;
    if (arc_index == 1496) return "W"  ;
    if (arc_index == 1497) return "E"  ;
    if (arc_index == 1498) return "E"  ;
    if (arc_index == 1499) return "E"  ;
    if (arc_index == 1500) return "E"  ;
    if (arc_index == 1501) return "E"  ;
    if (arc_index == 1502) return "E"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1504) return "W"  ;
    if (arc_index == 1505) return "E"  ;
    if (arc_index == 1506) return "E"  ;
    if (arc_index == 1507) return "E"  ;
    if (arc_index == 1508) return "E"  ;
    if (arc_index == 1509) return "E"  ;
    if (arc_index == 1510) return "E"  ;
    if (arc_index == 1511) return "E"  ;
    if (arc_index == 1512) return "E"  ;
    if (arc_index == 1513) return "E"  ;
    if (arc_index == 1514) return "E"  ;
    if (arc_index == 1515) return "E"  ;
    if (arc_index == 1516) return "W"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1529) return "H"  ;
    if (arc_index == 1546) return "H"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1574) return "H"  ;
    if (arc_index == 1592) return "H"  ;
    if (arc_index == 1710) return "H"  ;
    if (arc_index == 1723) return "E"  ;
    if (arc_index == 1773) return "H"  ;
    if (arc_index == 1810) return "H"  ;
    if (arc_index == 1855) return "H"  ;
    if (arc_index == 1950) return "H"  ;
    if (arc_index == 2017) return "E"  ;
    if (arc_index == 2018) return "E"  ;
    if (arc_index == 2019) return "E"  ;
    if (arc_index == 2034) return "H"  ;
    if (arc_index == 2080) return "H"  ;
    if (arc_index == 2119) return "E"  ;
    if (arc_index == 2143) return "H"  ;
    if (arc_index == 2150) return "E"  ;
    if (arc_index == 2151) return "E"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2180) return "W"  ;
    if (arc_index == 2212) return "W"  ;
    if (arc_index == 2259) return "H"  ;
    if (arc_index == 2348) return "H"  ;
    if (arc_index == 2350) return "H"  ;
    if (arc_index == 2362) return "H"  ;
    if (arc_index == 2377) return "W"  ;
    if (arc_index == 2444) return "E"  ;
    if (arc_index == 2446) return "E"  ;
    if (arc_index == 2447) return "E"  ;
    if (arc_index == 2448) return "E"  ;
    if (arc_index == 2449) return "E"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2455) return "E"  ;
    if (arc_index == 2462) return "E"  ;
    if (arc_index == 2483) return "E"  ;
    if (arc_index == 2491) return "E"  ;
    if (arc_index == 2493) return "H"  ;
    if (arc_index == 2513) return "E"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2577) return "E"  ;
    if (arc_index == 2578) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2646) return "H"  ;
    if (arc_index == 2704) return "H"  ;
    if (arc_index == 2815) return "H"  ;
    if (arc_index == 2885) return "H"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 0)) begin 
    if (arc_index == 135) return "H"  ;
    if (arc_index == 383) return "H"  ;
    if (arc_index == 391) return "H"  ;
    if (arc_index == 487) return "E"  ;
    if (arc_index == 491) return "E"  ;
    if (arc_index == 500) return "E"  ;
    if (arc_index == 505) return "E"  ;
    if (arc_index == 546) return "H"  ;
    if (arc_index == 575) return "E"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 679) return "H"  ;
    if (arc_index == 687) return "H"  ;
    if (arc_index == 774) return "H"  ;
    if (arc_index == 900) return "H"  ;
    if (arc_index == 947) return "H"  ;
    if (arc_index == 1011) return "H"  ;
    if (arc_index == 1022) return "H"  ;
    if (arc_index == 1081) return "H"  ;
    if (arc_index == 1256) return "H"  ;
    if (arc_index == 1453) return "H"  ;
    if (arc_index == 1496) return "H"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1519) return "E"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1522) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1524) return "E"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1526) return "E"  ;
    if (arc_index == 1527) return "E"  ;
    if (arc_index == 1528) return "E"  ;
    if (arc_index == 1529) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1532) return "E"  ;
    if (arc_index == 1533) return "E"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1535) return "E"  ;
    if (arc_index == 1536) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1538) return "E"  ;
    if (arc_index == 1539) return "E"  ;
    if (arc_index == 1551) return "H"  ;
    if (arc_index == 1562) return "H"  ;
    if (arc_index == 1589) return "E"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1596) return "H"  ;
    if (arc_index == 1602) return "E"  ;
    if (arc_index == 1603) return "E"  ;
    if (arc_index == 1795) return "H"  ;
    if (arc_index == 1972) return "H"  ;
    if (arc_index == 2056) return "H"  ;
    if (arc_index == 2165) return "H"  ;
    if (arc_index == 2281) return "H"  ;
    if (arc_index == 2370) return "H"  ;
    if (arc_index == 2384) return "H"  ;
    if (arc_index == 2436) return "H"  ;
    if (arc_index == 2515) return "H"  ;
    if (arc_index == 2581) return "H"  ;
    if (arc_index == 2668) return "H"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 11)) begin 
    if (arc_index == 146) return "H"  ;
    if (arc_index == 168) return "H"  ;
    if (arc_index == 230) return "H"  ;
    if (arc_index == 318) return "H"  ;
    if (arc_index == 413) return "H"  ;
    if (arc_index == 447) return "H"  ;
    if (arc_index == 544) return "H"  ;
    if (arc_index == 566) return "H"  ;
    if (arc_index == 568) return "H"  ;
    if (arc_index == 597) return "H"  ;
    if (arc_index == 630) return "W"  ;
    if (arc_index == 632) return "W"  ;
    if (arc_index == 701) return "H"  ;
    if (arc_index == 709) return "H"  ;
    if (arc_index == 711) return "H"  ;
    if (arc_index == 796) return "H"  ;
    if (arc_index == 922) return "H"  ;
    if (arc_index == 1033) return "H"  ;
    if (arc_index == 1034) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1048) return "W"  ;
    if (arc_index == 1049) return "W"  ;
    if (arc_index == 1050) return "W"  ;
    if (arc_index == 1103) return "H"  ;
    if (arc_index == 1128) return "H"  ;
    if (arc_index == 1249) return "H"  ;
    if (arc_index == 1278) return "H"  ;
    if (arc_index == 1475) return "H"  ;
    if (arc_index == 1518) return "H"  ;
    if (arc_index == 1537) return "H"  ;
    if (arc_index == 1540) return "H"  ;
    if (arc_index == 1541) return "W"  ;
    if (arc_index == 1542) return "W"  ;
    if (arc_index == 1543) return "W"  ;
    if (arc_index == 1544) return "W"  ;
    if (arc_index == 1545) return "W"  ;
    if (arc_index == 1546) return "W"  ;
    if (arc_index == 1547) return "W"  ;
    if (arc_index == 1548) return "W"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1552) return "W"  ;
    if (arc_index == 1553) return "W"  ;
    if (arc_index == 1554) return "W"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1556) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1558) return "W"  ;
    if (arc_index == 1559) return "W"  ;
    if (arc_index == 1560) return "W"  ;
    if (arc_index == 1561) return "W"  ;
    if (arc_index == 1573) return "H"  ;
    if (arc_index == 1618) return "H"  ;
    if (arc_index == 1817) return "H"  ;
    if (arc_index == 1874) return "H"  ;
    if (arc_index == 1994) return "H"  ;
    if (arc_index == 2073) return "H"  ;
    if (arc_index == 2078) return "H"  ;
    if (arc_index == 2114) return "H"  ;
    if (arc_index == 2187) return "H"  ;
    if (arc_index == 2303) return "H"  ;
    if (arc_index == 2311) return "H"  ;
    if (arc_index == 2378) return "H"  ;
    if (arc_index == 2388) return "H"  ;
    if (arc_index == 2392) return "H"  ;
    if (arc_index == 2396) return "H"  ;
    if (arc_index == 2406) return "H"  ;
    if (arc_index == 2409) return "H"  ;
    if (arc_index == 2537) return "H"  ;
    if (arc_index == 2618) return "H"  ;
    if (arc_index == 2621) return "H"  ;
    if (arc_index == 2642) return "H"  ;
    if (arc_index == 2651) return "H"  ;
    if (arc_index == 2653) return "H"  ;
    if (arc_index == 2658) return "H"  ;
    if (arc_index == 2690) return "H"  ;
    if (arc_index == 2711) return "H"  ;
    if (arc_index == 2724) return "H"  ;
    if (arc_index == 2727) return "H"  ;
    if (arc_index == 2833) return "H"  ;
    if (arc_index == 2908) return "W"  ;
    if (arc_index == 2917) return "W"  ;
    if (arc_index == 2921) return "W"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 10)) begin 
    if (arc_index == 252) return "E"  ;
    if (arc_index == 361) return "E"  ;
    if (arc_index == 435) return "H"  ;
    if (arc_index == 590) return "H"  ;
    if (arc_index == 723) return "H"  ;
    if (arc_index == 731) return "H"  ;
    if (arc_index == 818) return "H"  ;
    if (arc_index == 864) return "E"  ;
    if (arc_index == 944) return "H"  ;
    if (arc_index == 1055) return "H"  ;
    if (arc_index == 1125) return "H"  ;
    if (arc_index == 1300) return "H"  ;
    if (arc_index == 1497) return "H"  ;
    if (arc_index == 1513) return "E"  ;
    if (arc_index == 1540) return "H"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1565) return "W"  ;
    if (arc_index == 1566) return "W"  ;
    if (arc_index == 1567) return "W"  ;
    if (arc_index == 1568) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1570) return "W"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1572) return "W"  ;
    if (arc_index == 1573) return "W"  ;
    if (arc_index == 1574) return "W"  ;
    if (arc_index == 1575) return "W"  ;
    if (arc_index == 1576) return "W"  ;
    if (arc_index == 1577) return "W"  ;
    if (arc_index == 1578) return "W"  ;
    if (arc_index == 1579) return "W"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1581) return "W"  ;
    if (arc_index == 1582) return "W"  ;
    if (arc_index == 1583) return "W"  ;
    if (arc_index == 1595) return "H"  ;
    if (arc_index == 1640) return "H"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1839) return "H"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2016) return "H"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2100) return "H"  ;
    if (arc_index == 2209) return "H"  ;
    if (arc_index == 2325) return "H"  ;
    if (arc_index == 2414) return "H"  ;
    if (arc_index == 2428) return "H"  ;
    if (arc_index == 2559) return "H"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2646) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2657) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2660) return "W"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2712) return "H"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 0)) begin 
    if (arc_index == 135) return "H"  ;
    if (arc_index == 388) return "H"  ;
    if (arc_index == 457) return "H"  ;
    if (arc_index == 485) return "H"  ;
    if (arc_index == 486) return "E"  ;
    if (arc_index == 492) return "E"  ;
    if (arc_index == 493) return "E"  ;
    if (arc_index == 494) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 575) return "E"  ;
    if (arc_index == 579) return "E"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 582) return "E"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 588) return "E"  ;
    if (arc_index == 592) return "E"  ;
    if (arc_index == 612) return "H"  ;
    if (arc_index == 745) return "H"  ;
    if (arc_index == 753) return "H"  ;
    if (arc_index == 761) return "H"  ;
    if (arc_index == 840) return "H"  ;
    if (arc_index == 947) return "H"  ;
    if (arc_index == 957) return "H"  ;
    if (arc_index == 966) return "H"  ;
    if (arc_index == 1026) return "H"  ;
    if (arc_index == 1077) return "H"  ;
    if (arc_index == 1081) return "H"  ;
    if (arc_index == 1147) return "H"  ;
    if (arc_index == 1219) return "H"  ;
    if (arc_index == 1322) return "H"  ;
    if (arc_index == 1453) return "H"  ;
    if (arc_index == 1481) return "H"  ;
    if (arc_index == 1519) return "H"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1562) return "H"  ;
    if (arc_index == 1584) return "E"  ;
    if (arc_index == 1585) return "E"  ;
    if (arc_index == 1586) return "E"  ;
    if (arc_index == 1587) return "E"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1589) return "E"  ;
    if (arc_index == 1590) return "E"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1593) return "E"  ;
    if (arc_index == 1594) return "E"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1596) return "E"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1599) return "E"  ;
    if (arc_index == 1600) return "E"  ;
    if (arc_index == 1601) return "E"  ;
    if (arc_index == 1602) return "E"  ;
    if (arc_index == 1603) return "E"  ;
    if (arc_index == 1604) return "E"  ;
    if (arc_index == 1605) return "E"  ;
    if (arc_index == 1617) return "H"  ;
    if (arc_index == 1662) return "H"  ;
    if (arc_index == 1861) return "H"  ;
    if (arc_index == 1918) return "H"  ;
    if (arc_index == 2021) return "H"  ;
    if (arc_index == 2038) return "H"  ;
    if (arc_index == 2044) return "H"  ;
    if (arc_index == 2122) return "H"  ;
    if (arc_index == 2231) return "H"  ;
    if (arc_index == 2347) return "H"  ;
    if (arc_index == 2423) return "H"  ;
    if (arc_index == 2436) return "H"  ;
    if (arc_index == 2450) return "H"  ;
    if (arc_index == 2571) return "H"  ;
    if (arc_index == 2581) return "H"  ;
    if (arc_index == 2663) return "H"  ;
    if (arc_index == 2667) return "H"  ;
    if (arc_index == 2671) return "H"  ;
    if (arc_index == 2674) return "H"  ;
    if (arc_index == 2678) return "H"  ;
    if (arc_index == 2679) return "H"  ;
    if (arc_index == 2695) return "H"  ;
    if (arc_index == 2734) return "H"  ;
    if (arc_index == 2740) return "H"  ;
    if (arc_index == 2792) return "H"  ;
    if (arc_index == 2863) return "E"  ;
    if (arc_index == 2874) return "E"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2879) return "E"  ;
    if (arc_index == 2903) return "E"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 4)) begin 
    if (arc_index == 26) return "E"  ;
    if (arc_index == 28) return "E"  ;
    if (arc_index == 51) return "E"  ;
    if (arc_index == 58) return "E"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 86) return "E"  ;
    if (arc_index == 101) return "E"  ;
    if (arc_index == 123) return "E"  ;
    if (arc_index == 136) return "W"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 362) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 442) return "W"  ;
    if (arc_index == 456) return "W"  ;
    if (arc_index == 475) return "E"  ;
    if (arc_index == 479) return "H"  ;
    if (arc_index == 480) return "E"  ;
    if (arc_index == 482) return "E"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 512) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 535) return "E"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 593) return "E"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 609) return "W"  ;
    if (arc_index == 634) return "H"  ;
    if (arc_index == 676) return "H"  ;
    if (arc_index == 693) return "H"  ;
    if (arc_index == 717) return "H"  ;
    if (arc_index == 719) return "H"  ;
    if (arc_index == 726) return "H"  ;
    if (arc_index == 744) return "H"  ;
    if (arc_index == 752) return "H"  ;
    if (arc_index == 759) return "E"  ;
    if (arc_index == 767) return "H"  ;
    if (arc_index == 769) return "H"  ;
    if (arc_index == 775) return "H"  ;
    if (arc_index == 777) return "H"  ;
    if (arc_index == 819) return "W"  ;
    if (arc_index == 822) return "W"  ;
    if (arc_index == 862) return "H"  ;
    if (arc_index == 882) return "E"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 965) return "E"  ;
    if (arc_index == 972) return "E"  ;
    if (arc_index == 974) return "E"  ;
    if (arc_index == 988) return "H"  ;
    if (arc_index == 996) return "H"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1008) return "E"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1047) return "E"  ;
    if (arc_index == 1056) return "W"  ;
    if (arc_index == 1078) return "E"  ;
    if (arc_index == 1085) return "E"  ;
    if (arc_index == 1092) return "E"  ;
    if (arc_index == 1099) return "H"  ;
    if (arc_index == 1105) return "W"  ;
    if (arc_index == 1110) return "W"  ;
    if (arc_index == 1111) return "W"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1169) return "H"  ;
    if (arc_index == 1185) return "H"  ;
    if (arc_index == 1190) return "E"  ;
    if (arc_index == 1197) return "E"  ;
    if (arc_index == 1280) return "E"  ;
    if (arc_index == 1308) return "E"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1344) return "H"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1388) return "W"  ;
    if (arc_index == 1390) return "W"  ;
    if (arc_index == 1391) return "W"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1428) return "W"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1453) return "W"  ;
    if (arc_index == 1459) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1541) return "H"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1584) return "H"  ;
    if (arc_index == 1586) return "E"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1606) return "E"  ;
    if (arc_index == 1607) return "E"  ;
    if (arc_index == 1608) return "E"  ;
    if (arc_index == 1609) return "E"  ;
    if (arc_index == 1610) return "E"  ;
    if (arc_index == 1611) return "E"  ;
    if (arc_index == 1612) return "W"  ;
    if (arc_index == 1613) return "E"  ;
    if (arc_index == 1614) return "E"  ;
    if (arc_index == 1615) return "E"  ;
    if (arc_index == 1616) return "W"  ;
    if (arc_index == 1617) return "W"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1619) return "E"  ;
    if (arc_index == 1620) return "E"  ;
    if (arc_index == 1621) return "E"  ;
    if (arc_index == 1622) return "W"  ;
    if (arc_index == 1623) return "W"  ;
    if (arc_index == 1624) return "E"  ;
    if (arc_index == 1625) return "E"  ;
    if (arc_index == 1626) return "E"  ;
    if (arc_index == 1627) return "E"  ;
    if (arc_index == 1638) return "E"  ;
    if (arc_index == 1639) return "H"  ;
    if (arc_index == 1645) return "H"  ;
    if (arc_index == 1650) return "E"  ;
    if (arc_index == 1653) return "E"  ;
    if (arc_index == 1654) return "E"  ;
    if (arc_index == 1655) return "E"  ;
    if (arc_index == 1663) return "E"  ;
    if (arc_index == 1666) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1670) return "E"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1673) return "W"  ;
    if (arc_index == 1684) return "H"  ;
    if (arc_index == 1697) return "H"  ;
    if (arc_index == 1741) return "H"  ;
    if (arc_index == 1747) return "E"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1755) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1784) return "E"  ;
    if (arc_index == 1790) return "W"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1804) return "W"  ;
    if (arc_index == 1822) return "W"  ;
    if (arc_index == 1829) return "E"  ;
    if (arc_index == 1849) return "W"  ;
    if (arc_index == 1853) return "W"  ;
    if (arc_index == 1857) return "W"  ;
    if (arc_index == 1861) return "W"  ;
    if (arc_index == 1883) return "H"  ;
    if (arc_index == 1892) return "W"  ;
    if (arc_index == 1898) return "W"  ;
    if (arc_index == 1904) return "W"  ;
    if (arc_index == 1911) return "W"  ;
    if (arc_index == 1916) return "W"  ;
    if (arc_index == 1917) return "E"  ;
    if (arc_index == 1922) return "E"  ;
    if (arc_index == 1924) return "E"  ;
    if (arc_index == 1925) return "E"  ;
    if (arc_index == 1926) return "E"  ;
    if (arc_index == 1928) return "E"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1946) return "E"  ;
    if (arc_index == 1952) return "E"  ;
    if (arc_index == 1980) return "E"  ;
    if (arc_index == 1981) return "E"  ;
    if (arc_index == 1983) return "E"  ;
    if (arc_index == 1994) return "E"  ;
    if (arc_index == 1998) return "E"  ;
    if (arc_index == 2006) return "E"  ;
    if (arc_index == 2013) return "E"  ;
    if (arc_index == 2023) return "E"  ;
    if (arc_index == 2032) return "E"  ;
    if (arc_index == 2036) return "E"  ;
    if (arc_index == 2042) return "E"  ;
    if (arc_index == 2050) return "E"  ;
    if (arc_index == 2055) return "E"  ;
    if (arc_index == 2057) return "E"  ;
    if (arc_index == 2058) return "E"  ;
    if (arc_index == 2060) return "H"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2104) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2115) return "W"  ;
    if (arc_index == 2132) return "W"  ;
    if (arc_index == 2144) return "H"  ;
    if (arc_index == 2148) return "H"  ;
    if (arc_index == 2149) return "H"  ;
    if (arc_index == 2152) return "E"  ;
    if (arc_index == 2154) return "E"  ;
    if (arc_index == 2188) return "W"  ;
    if (arc_index == 2202) return "W"  ;
    if (arc_index == 2223) return "W"  ;
    if (arc_index == 2224) return "E"  ;
    if (arc_index == 2236) return "E"  ;
    if (arc_index == 2238) return "E"  ;
    if (arc_index == 2243) return "E"  ;
    if (arc_index == 2253) return "H"  ;
    if (arc_index == 2254) return "H"  ;
    if (arc_index == 2276) return "H"  ;
    if (arc_index == 2280) return "W"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2313) return "W"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2363) return "W"  ;
    if (arc_index == 2368) return "W"  ;
    if (arc_index == 2369) return "H"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2375) return "W"  ;
    if (arc_index == 2413) return "W"  ;
    if (arc_index == 2457) return "W"  ;
    if (arc_index == 2458) return "H"  ;
    if (arc_index == 2472) return "H"  ;
    if (arc_index == 2486) return "H"  ;
    if (arc_index == 2494) return "W"  ;
    if (arc_index == 2499) return "W"  ;
    if (arc_index == 2502) return "W"  ;
    if (arc_index == 2508) return "W"  ;
    if (arc_index == 2510) return "W"  ;
    if (arc_index == 2518) return "W"  ;
    if (arc_index == 2519) return "E"  ;
    if (arc_index == 2540) return "W"  ;
    if (arc_index == 2574) return "W"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2603) return "H"  ;
    if (arc_index == 2607) return "H"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2685) return "W"  ;
    if (arc_index == 2691) return "W"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2706) return "E"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2752) return "E"  ;
    if (arc_index == 2754) return "W"  ;
    if (arc_index == 2755) return "W"  ;
    if (arc_index == 2756) return "H"  ;
    if (arc_index == 2758) return "E"  ;
    if (arc_index == 2759) return "E"  ;
    if (arc_index == 2762) return "W"  ;
    if (arc_index == 2764) return "E"  ;
    if (arc_index == 2766) return "W"  ;
    if (arc_index == 2767) return "E"  ;
    if (arc_index == 2771) return "E"  ;
    if (arc_index == 2774) return "E"  ;
    if (arc_index == 2778) return "W"  ;
    if (arc_index == 2781) return "W"  ;
    if (arc_index == 2785) return "W"  ;
    if (arc_index == 2789) return "W"  ;
    if (arc_index == 2793) return "W"  ;
    if (arc_index == 2801) return "E"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2809) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2817) return "E"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2882) return "E"  ;
    if (arc_index == 2888) return "E"  ;
    if (arc_index == 2890) return "E"  ;
    if (arc_index == 2892) return "E"  ;
    if (arc_index == 2893) return "E"  ;
    if (arc_index == 2899) return "E"  ;
    if (arc_index == 2900) return "W"  ;
    if (arc_index == 2901) return "W"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 2)) begin 
    if (arc_index == 7) return "W"  ;
    if (arc_index == 65) return "W"  ;
    if (arc_index == 76) return "E"  ;
    if (arc_index == 79) return "W"  ;
    if (arc_index == 80) return "W"  ;
    if (arc_index == 106) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 115) return "W"  ;
    if (arc_index == 138) return "W"  ;
    if (arc_index == 160) return "W"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 384) return "W"  ;
    if (arc_index == 390) return "W"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 443) return "E"  ;
    if (arc_index == 494) return "E"  ;
    if (arc_index == 501) return "H"  ;
    if (arc_index == 503) return "H"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 520) return "E"  ;
    if (arc_index == 521) return "E"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 591) return "E"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 654) return "W"  ;
    if (arc_index == 656) return "H"  ;
    if (arc_index == 668) return "H"  ;
    if (arc_index == 717) return "H"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 751) return "W"  ;
    if (arc_index == 770) return "W"  ;
    if (arc_index == 779) return "W"  ;
    if (arc_index == 789) return "H"  ;
    if (arc_index == 797) return "H"  ;
    if (arc_index == 799) return "H"  ;
    if (arc_index == 803) return "H"  ;
    if (arc_index == 808) return "E"  ;
    if (arc_index == 858) return "E"  ;
    if (arc_index == 865) return "E"  ;
    if (arc_index == 877) return "E"  ;
    if (arc_index == 880) return "E"  ;
    if (arc_index == 884) return "H"  ;
    if (arc_index == 886) return "H"  ;
    if (arc_index == 888) return "E"  ;
    if (arc_index == 896) return "E"  ;
    if (arc_index == 900) return "E"  ;
    if (arc_index == 906) return "E"  ;
    if (arc_index == 907) return "E"  ;
    if (arc_index == 908) return "E"  ;
    if (arc_index == 909) return "E"  ;
    if (arc_index == 913) return "E"  ;
    if (arc_index == 931) return "E"  ;
    if (arc_index == 942) return "E"  ;
    if (arc_index == 946) return "E"  ;
    if (arc_index == 953) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 1010) return "H"  ;
    if (arc_index == 1075) return "H"  ;
    if (arc_index == 1077) return "W"  ;
    if (arc_index == 1105) return "W"  ;
    if (arc_index == 1121) return "H"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1170) return "W"  ;
    if (arc_index == 1191) return "H"  ;
    if (arc_index == 1192) return "W"  ;
    if (arc_index == 1193) return "W"  ;
    if (arc_index == 1202) return "W"  ;
    if (arc_index == 1208) return "E"  ;
    if (arc_index == 1209) return "E"  ;
    if (arc_index == 1213) return "E"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1231) return "E"  ;
    if (arc_index == 1296) return "E"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1366) return "H"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1438) return "W"  ;
    if (arc_index == 1465) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1527) return "W"  ;
    if (arc_index == 1533) return "W"  ;
    if (arc_index == 1563) return "H"  ;
    if (arc_index == 1569) return "H"  ;
    if (arc_index == 1584) return "H"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1594) return "E"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1599) return "E"  ;
    if (arc_index == 1605) return "E"  ;
    if (arc_index == 1606) return "H"  ;
    if (arc_index == 1617) return "W"  ;
    if (arc_index == 1628) return "W"  ;
    if (arc_index == 1629) return "E"  ;
    if (arc_index == 1630) return "E"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1633) return "E"  ;
    if (arc_index == 1634) return "E"  ;
    if (arc_index == 1635) return "E"  ;
    if (arc_index == 1636) return "E"  ;
    if (arc_index == 1637) return "E"  ;
    if (arc_index == 1638) return "E"  ;
    if (arc_index == 1639) return "E"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1641) return "E"  ;
    if (arc_index == 1642) return "E"  ;
    if (arc_index == 1643) return "E"  ;
    if (arc_index == 1644) return "E"  ;
    if (arc_index == 1645) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1647) return "E"  ;
    if (arc_index == 1648) return "E"  ;
    if (arc_index == 1649) return "E"  ;
    if (arc_index == 1661) return "H"  ;
    if (arc_index == 1664) return "H"  ;
    if (arc_index == 1665) return "H"  ;
    if (arc_index == 1674) return "W"  ;
    if (arc_index == 1706) return "H"  ;
    if (arc_index == 1719) return "H"  ;
    if (arc_index == 1723) return "H"  ;
    if (arc_index == 1726) return "H"  ;
    if (arc_index == 1731) return "E"  ;
    if (arc_index == 1735) return "E"  ;
    if (arc_index == 1740) return "E"  ;
    if (arc_index == 1743) return "E"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1754) return "E"  ;
    if (arc_index == 1768) return "E"  ;
    if (arc_index == 1830) return "W"  ;
    if (arc_index == 1831) return "W"  ;
    if (arc_index == 1835) return "W"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1897) return "W"  ;
    if (arc_index == 1905) return "H"  ;
    if (arc_index == 1914) return "W"  ;
    if (arc_index == 1921) return "W"  ;
    if (arc_index == 1923) return "E"  ;
    if (arc_index == 1929) return "E"  ;
    if (arc_index == 1931) return "E"  ;
    if (arc_index == 1935) return "E"  ;
    if (arc_index == 1936) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1940) return "E"  ;
    if (arc_index == 1946) return "E"  ;
    if (arc_index == 1947) return "E"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1949) return "E"  ;
    if (arc_index == 1952) return "E"  ;
    if (arc_index == 1953) return "E"  ;
    if (arc_index == 1954) return "E"  ;
    if (arc_index == 1969) return "W"  ;
    if (arc_index == 2002) return "W"  ;
    if (arc_index == 2007) return "W"  ;
    if (arc_index == 2015) return "W"  ;
    if (arc_index == 2082) return "H"  ;
    if (arc_index == 2122) return "W"  ;
    if (arc_index == 2166) return "H"  ;
    if (arc_index == 2191) return "H"  ;
    if (arc_index == 2223) return "H"  ;
    if (arc_index == 2224) return "E"  ;
    if (arc_index == 2238) return "E"  ;
    if (arc_index == 2275) return "H"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "H"  ;
    if (arc_index == 2452) return "H"  ;
    if (arc_index == 2469) return "H"  ;
    if (arc_index == 2480) return "H"  ;
    if (arc_index == 2494) return "H"  ;
    if (arc_index == 2526) return "H"  ;
    if (arc_index == 2555) return "H"  ;
    if (arc_index == 2566) return "E"  ;
    if (arc_index == 2576) return "E"  ;
    if (arc_index == 2582) return "E"  ;
    if (arc_index == 2590) return "E"  ;
    if (arc_index == 2597) return "E"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2625) return "H"  ;
    if (arc_index == 2670) return "E"  ;
    if (arc_index == 2677) return "E"  ;
    if (arc_index == 2688) return "E"  ;
    if (arc_index == 2695) return "W"  ;
    if (arc_index == 2699) return "W"  ;
    if (arc_index == 2701) return "W"  ;
    if (arc_index == 2733) return "W"  ;
    if (arc_index == 2746) return "W"  ;
    if (arc_index == 2765) return "W"  ;
    if (arc_index == 2778) return "H"  ;
    if (arc_index == 2788) return "W"  ;
    if (arc_index == 2812) return "W"  ;
    if (arc_index == 2860) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2868) return "E"  ;
    if (arc_index == 2903) return "W"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 3)) begin 
    if (arc_index == 41) return "W"  ;
    if (arc_index == 49) return "W"  ;
    if (arc_index == 50) return "W"  ;
    if (arc_index == 76) return "W"  ;
    if (arc_index == 136) return "W"  ;
    if (arc_index == 152) return "W"  ;
    if (arc_index == 200) return "W"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 384) return "W"  ;
    if (arc_index == 390) return "W"  ;
    if (arc_index == 404) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 470) return "W"  ;
    if (arc_index == 471) return "W"  ;
    if (arc_index == 472) return "W"  ;
    if (arc_index == 478) return "W"  ;
    if (arc_index == 479) return "E"  ;
    if (arc_index == 480) return "E"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 512) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 523) return "H"  ;
    if (arc_index == 525) return "H"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 572) return "W"  ;
    if (arc_index == 574) return "W"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 593) return "E"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 664) return "W"  ;
    if (arc_index == 675) return "W"  ;
    if (arc_index == 678) return "H"  ;
    if (arc_index == 750) return "H"  ;
    if (arc_index == 755) return "H"  ;
    if (arc_index == 785) return "H"  ;
    if (arc_index == 810) return "H"  ;
    if (arc_index == 811) return "H"  ;
    if (arc_index == 819) return "H"  ;
    if (arc_index == 890) return "H"  ;
    if (arc_index == 895) return "H"  ;
    if (arc_index == 898) return "H"  ;
    if (arc_index == 906) return "H"  ;
    if (arc_index == 909) return "H"  ;
    if (arc_index == 914) return "H"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 965) return "E"  ;
    if (arc_index == 987) return "E"  ;
    if (arc_index == 994) return "W"  ;
    if (arc_index == 995) return "W"  ;
    if (arc_index == 1032) return "H"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1056) return "W"  ;
    if (arc_index == 1085) return "E"  ;
    if (arc_index == 1092) return "E"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1099) return "E"  ;
    if (arc_index == 1105) return "W"  ;
    if (arc_index == 1110) return "W"  ;
    if (arc_index == 1111) return "W"  ;
    if (arc_index == 1143) return "H"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1208) return "W"  ;
    if (arc_index == 1213) return "H"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1279) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1388) return "H"  ;
    if (arc_index == 1391) return "W"  ;
    if (arc_index == 1407) return "W"  ;
    if (arc_index == 1453) return "W"  ;
    if (arc_index == 1465) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1477) return "W"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1564) return "E"  ;
    if (arc_index == 1584) return "E"  ;
    if (arc_index == 1585) return "H"  ;
    if (arc_index == 1586) return "E"  ;
    if (arc_index == 1587) return "E"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1599) return "E"  ;
    if (arc_index == 1612) return "E"  ;
    if (arc_index == 1616) return "W"  ;
    if (arc_index == 1622) return "W"  ;
    if (arc_index == 1628) return "H"  ;
    if (arc_index == 1629) return "H"  ;
    if (arc_index == 1633) return "H"  ;
    if (arc_index == 1639) return "E"  ;
    if (arc_index == 1650) return "E"  ;
    if (arc_index == 1651) return "E"  ;
    if (arc_index == 1652) return "W"  ;
    if (arc_index == 1653) return "E"  ;
    if (arc_index == 1654) return "E"  ;
    if (arc_index == 1655) return "E"  ;
    if (arc_index == 1656) return "W"  ;
    if (arc_index == 1657) return "W"  ;
    if (arc_index == 1658) return "W"  ;
    if (arc_index == 1659) return "W"  ;
    if (arc_index == 1660) return "W"  ;
    if (arc_index == 1661) return "W"  ;
    if (arc_index == 1662) return "W"  ;
    if (arc_index == 1663) return "E"  ;
    if (arc_index == 1664) return "W"  ;
    if (arc_index == 1665) return "W"  ;
    if (arc_index == 1666) return "E"  ;
    if (arc_index == 1667) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1669) return "E"  ;
    if (arc_index == 1670) return "E"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1673) return "W"  ;
    if (arc_index == 1683) return "H"  ;
    if (arc_index == 1712) return "H"  ;
    if (arc_index == 1715) return "H"  ;
    if (arc_index == 1724) return "H"  ;
    if (arc_index == 1728) return "H"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1753) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1790) return "E"  ;
    if (arc_index == 1804) return "E"  ;
    if (arc_index == 1822) return "E"  ;
    if (arc_index == 1827) return "E"  ;
    if (arc_index == 1829) return "E"  ;
    if (arc_index == 1830) return "W"  ;
    if (arc_index == 1831) return "W"  ;
    if (arc_index == 1834) return "W"  ;
    if (arc_index == 1835) return "W"  ;
    if (arc_index == 1839) return "W"  ;
    if (arc_index == 1842) return "W"  ;
    if (arc_index == 1843) return "W"  ;
    if (arc_index == 1845) return "W"  ;
    if (arc_index == 1849) return "W"  ;
    if (arc_index == 1853) return "W"  ;
    if (arc_index == 1861) return "W"  ;
    if (arc_index == 1892) return "W"  ;
    if (arc_index == 1916) return "E"  ;
    if (arc_index == 1917) return "E"  ;
    if (arc_index == 1922) return "E"  ;
    if (arc_index == 1924) return "E"  ;
    if (arc_index == 1925) return "E"  ;
    if (arc_index == 1926) return "E"  ;
    if (arc_index == 1927) return "H"  ;
    if (arc_index == 1928) return "E"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1941) return "E"  ;
    if (arc_index == 1987) return "E"  ;
    if (arc_index == 1992) return "W"  ;
    if (arc_index == 2001) return "W"  ;
    if (arc_index == 2007) return "W"  ;
    if (arc_index == 2023) return "E"  ;
    if (arc_index == 2024) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2035) return "E"  ;
    if (arc_index == 2036) return "E"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2040) return "E"  ;
    if (arc_index == 2042) return "E"  ;
    if (arc_index == 2043) return "E"  ;
    if (arc_index == 2075) return "E"  ;
    if (arc_index == 2104) return "H"  ;
    if (arc_index == 2115) return "W"  ;
    if (arc_index == 2170) return "W"  ;
    if (arc_index == 2171) return "W"  ;
    if (arc_index == 2188) return "H"  ;
    if (arc_index == 2202) return "H"  ;
    if (arc_index == 2223) return "E"  ;
    if (arc_index == 2238) return "E"  ;
    if (arc_index == 2280) return "E"  ;
    if (arc_index == 2297) return "H"  ;
    if (arc_index == 2363) return "H"  ;
    if (arc_index == 2368) return "W"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2413) return "H"  ;
    if (arc_index == 2434) return "H"  ;
    if (arc_index == 2442) return "H"  ;
    if (arc_index == 2460) return "W"  ;
    if (arc_index == 2469) return "W"  ;
    if (arc_index == 2475) return "W"  ;
    if (arc_index == 2477) return "W"  ;
    if (arc_index == 2483) return "W"  ;
    if (arc_index == 2485) return "W"  ;
    if (arc_index == 2494) return "W"  ;
    if (arc_index == 2499) return "W"  ;
    if (arc_index == 2502) return "H"  ;
    if (arc_index == 2516) return "H"  ;
    if (arc_index == 2540) return "H"  ;
    if (arc_index == 2557) return "H"  ;
    if (arc_index == 2589) return "H"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2647) return "H"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2678) return "W"  ;
    if (arc_index == 2692) return "W"  ;
    if (arc_index == 2702) return "W"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2754) return "W"  ;
    if (arc_index == 2762) return "W"  ;
    if (arc_index == 2766) return "W"  ;
    if (arc_index == 2770) return "W"  ;
    if (arc_index == 2778) return "W"  ;
    if (arc_index == 2793) return "W"  ;
    if (arc_index == 2800) return "H"  ;
    if (arc_index == 2801) return "E"  ;
    if (arc_index == 2803) return "E"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2809) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2842) return "E"  ;
    if (arc_index == 2854) return "E"  ;
    if (arc_index == 2856) return "E"  ;
    if (arc_index == 2861) return "E"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2881) return "E"  ;
    if (arc_index == 2900) return "W"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 8)) begin 
    if (arc_index == 24) return "E"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 89) return "E"  ;
    if (arc_index == 97) return "E"  ;
    if (arc_index == 109) return "E"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 154) return "E"  ;
    if (arc_index == 155) return "E"  ;
    if (arc_index == 163) return "E"  ;
    if (arc_index == 166) return "E"  ;
    if (arc_index == 171) return "E"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 183) return "W"  ;
    if (arc_index == 187) return "W"  ;
    if (arc_index == 198) return "W"  ;
    if (arc_index == 209) return "E"  ;
    if (arc_index == 219) return "E"  ;
    if (arc_index == 220) return "E"  ;
    if (arc_index == 225) return "E"  ;
    if (arc_index == 228) return "E"  ;
    if (arc_index == 230) return "E"  ;
    if (arc_index == 231) return "E"  ;
    if (arc_index == 232) return "E"  ;
    if (arc_index == 233) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 249) return "W"  ;
    if (arc_index == 250) return "E"  ;
    if (arc_index == 252) return "E"  ;
    if (arc_index == 253) return "E"  ;
    if (arc_index == 260) return "E"  ;
    if (arc_index == 271) return "E"  ;
    if (arc_index == 279) return "E"  ;
    if (arc_index == 282) return "E"  ;
    if (arc_index == 283) return "E"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 296) return "W"  ;
    if (arc_index == 297) return "W"  ;
    if (arc_index == 299) return "W"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 338) return "E"  ;
    if (arc_index == 339) return "E"  ;
    if (arc_index == 341) return "E"  ;
    if (arc_index == 420) return "E"  ;
    if (arc_index == 431) return "E"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 469) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 537) return "W"  ;
    if (arc_index == 538) return "W"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 541) return "W"  ;
    if (arc_index == 545) return "H"  ;
    if (arc_index == 547) return "H"  ;
    if (arc_index == 554) return "H"  ;
    if (arc_index == 599) return "H"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 660) return "W"  ;
    if (arc_index == 700) return "H"  ;
    if (arc_index == 704) return "H"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 730) return "W"  ;
    if (arc_index == 736) return "W"  ;
    if (arc_index == 758) return "W"  ;
    if (arc_index == 792) return "W"  ;
    if (arc_index == 801) return "W"  ;
    if (arc_index == 802) return "W"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 833) return "H"  ;
    if (arc_index == 841) return "H"  ;
    if (arc_index == 911) return "H"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 928) return "H"  ;
    if (arc_index == 929) return "H"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1040) return "E"  ;
    if (arc_index == 1052) return "E"  ;
    if (arc_index == 1054) return "H"  ;
    if (arc_index == 1073) return "H"  ;
    if (arc_index == 1086) return "H"  ;
    if (arc_index == 1130) return "H"  ;
    if (arc_index == 1134) return "H"  ;
    if (arc_index == 1136) return "H"  ;
    if (arc_index == 1140) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1165) return "H"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1235) return "H"  ;
    if (arc_index == 1236) return "H"  ;
    if (arc_index == 1239) return "H"  ;
    if (arc_index == 1255) return "E"  ;
    if (arc_index == 1257) return "E"  ;
    if (arc_index == 1259) return "E"  ;
    if (arc_index == 1261) return "E"  ;
    if (arc_index == 1263) return "E"  ;
    if (arc_index == 1274) return "W"  ;
    if (arc_index == 1275) return "W"  ;
    if (arc_index == 1277) return "E"  ;
    if (arc_index == 1304) return "E"  ;
    if (arc_index == 1313) return "W"  ;
    if (arc_index == 1332) return "W"  ;
    if (arc_index == 1340) return "W"  ;
    if (arc_index == 1354) return "W"  ;
    if (arc_index == 1363) return "W"  ;
    if (arc_index == 1410) return "H"  ;
    if (arc_index == 1436) return "E"  ;
    if (arc_index == 1474) return "E"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1488) return "E"  ;
    if (arc_index == 1489) return "E"  ;
    if (arc_index == 1501) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1541) return "W"  ;
    if (arc_index == 1542) return "W"  ;
    if (arc_index == 1543) return "W"  ;
    if (arc_index == 1546) return "W"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1553) return "W"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1595) return "W"  ;
    if (arc_index == 1607) return "H"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1650) return "H"  ;
    if (arc_index == 1668) return "H"  ;
    if (arc_index == 1671) return "H"  ;
    if (arc_index == 1672) return "H"  ;
    if (arc_index == 1673) return "H"  ;
    if (arc_index == 1674) return "W"  ;
    if (arc_index == 1675) return "W"  ;
    if (arc_index == 1676) return "W"  ;
    if (arc_index == 1677) return "W"  ;
    if (arc_index == 1678) return "W"  ;
    if (arc_index == 1679) return "W"  ;
    if (arc_index == 1680) return "W"  ;
    if (arc_index == 1681) return "E"  ;
    if (arc_index == 1682) return "E"  ;
    if (arc_index == 1683) return "W"  ;
    if (arc_index == 1684) return "W"  ;
    if (arc_index == 1685) return "W"  ;
    if (arc_index == 1686) return "W"  ;
    if (arc_index == 1687) return "W"  ;
    if (arc_index == 1688) return "W"  ;
    if (arc_index == 1689) return "W"  ;
    if (arc_index == 1690) return "W"  ;
    if (arc_index == 1691) return "W"  ;
    if (arc_index == 1692) return "W"  ;
    if (arc_index == 1693) return "W"  ;
    if (arc_index == 1705) return "H"  ;
    if (arc_index == 1708) return "H"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1750) return "H"  ;
    if (arc_index == 1763) return "H"  ;
    if (arc_index == 1792) return "H"  ;
    if (arc_index == 1805) return "H"  ;
    if (arc_index == 1809) return "H"  ;
    if (arc_index == 1836) return "H"  ;
    if (arc_index == 1867) return "H"  ;
    if (arc_index == 1870) return "W"  ;
    if (arc_index == 1874) return "E"  ;
    if (arc_index == 1882) return "E"  ;
    if (arc_index == 1888) return "E"  ;
    if (arc_index == 1901) return "E"  ;
    if (arc_index == 1903) return "E"  ;
    if (arc_index == 1949) return "H"  ;
    if (arc_index == 1961) return "E"  ;
    if (arc_index == 1962) return "E"  ;
    if (arc_index == 1964) return "E"  ;
    if (arc_index == 1967) return "E"  ;
    if (arc_index == 1974) return "E"  ;
    if (arc_index == 1975) return "E"  ;
    if (arc_index == 1994) return "E"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 2063) return "E"  ;
    if (arc_index == 2072) return "E"  ;
    if (arc_index == 2079) return "W"  ;
    if (arc_index == 2098) return "W"  ;
    if (arc_index == 2106) return "W"  ;
    if (arc_index == 2114) return "E"  ;
    if (arc_index == 2126) return "H"  ;
    if (arc_index == 2172) return "E"  ;
    if (arc_index == 2182) return "E"  ;
    if (arc_index == 2188) return "W"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2210) return "H"  ;
    if (arc_index == 2214) return "H"  ;
    if (arc_index == 2215) return "H"  ;
    if (arc_index == 2218) return "H"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2267) return "E"  ;
    if (arc_index == 2288) return "E"  ;
    if (arc_index == 2307) return "E"  ;
    if (arc_index == 2313) return "E"  ;
    if (arc_index == 2319) return "H"  ;
    if (arc_index == 2322) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2344) return "W"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2361) return "W"  ;
    if (arc_index == 2372) return "W"  ;
    if (arc_index == 2398) return "W"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2402) return "W"  ;
    if (arc_index == 2412) return "W"  ;
    if (arc_index == 2416) return "W"  ;
    if (arc_index == 2435) return "H"  ;
    if (arc_index == 2446) return "H"  ;
    if (arc_index == 2454) return "H"  ;
    if (arc_index == 2462) return "H"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2524) return "H"  ;
    if (arc_index == 2538) return "H"  ;
    if (arc_index == 2599) return "H"  ;
    if (arc_index == 2600) return "H"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2669) return "H"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2705) return "E"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2714) return "W"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2739) return "W"  ;
    if (arc_index == 2784) return "W"  ;
    if (arc_index == 2822) return "H"  ;
    if (arc_index == 2840) return "H"  ;
    if (arc_index == 2847) return "H"  ;
    if (arc_index == 2848) return "H"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2907) return "E"  ;
    if (arc_index == 2908) return "E"  ;
    if (arc_index == 2913) return "E"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 5)) begin 
    if (arc_index == 164) return "W"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 550) return "W"  ;
    if (arc_index == 555) return "W"  ;
    if (arc_index == 559) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 565) return "W"  ;
    if (arc_index == 567) return "H"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 571) return "W"  ;
    if (arc_index == 577) return "E"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 664) return "E"  ;
    if (arc_index == 698) return "W"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 712) return "W"  ;
    if (arc_index == 722) return "H"  ;
    if (arc_index == 788) return "E"  ;
    if (arc_index == 790) return "E"  ;
    if (arc_index == 855) return "H"  ;
    if (arc_index == 863) return "H"  ;
    if (arc_index == 950) return "H"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 1076) return "H"  ;
    if (arc_index == 1187) return "H"  ;
    if (arc_index == 1197) return "E"  ;
    if (arc_index == 1257) return "H"  ;
    if (arc_index == 1386) return "E"  ;
    if (arc_index == 1408) return "E"  ;
    if (arc_index == 1417) return "W"  ;
    if (arc_index == 1418) return "W"  ;
    if (arc_index == 1419) return "W"  ;
    if (arc_index == 1424) return "W"  ;
    if (arc_index == 1425) return "W"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1432) return "H"  ;
    if (arc_index == 1441) return "E"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1629) return "H"  ;
    if (arc_index == 1672) return "H"  ;
    if (arc_index == 1694) return "H"  ;
    if (arc_index == 1695) return "E"  ;
    if (arc_index == 1696) return "E"  ;
    if (arc_index == 1697) return "E"  ;
    if (arc_index == 1698) return "E"  ;
    if (arc_index == 1699) return "E"  ;
    if (arc_index == 1700) return "E"  ;
    if (arc_index == 1701) return "E"  ;
    if (arc_index == 1702) return "E"  ;
    if (arc_index == 1703) return "E"  ;
    if (arc_index == 1704) return "E"  ;
    if (arc_index == 1705) return "E"  ;
    if (arc_index == 1706) return "W"  ;
    if (arc_index == 1707) return "W"  ;
    if (arc_index == 1708) return "E"  ;
    if (arc_index == 1709) return "W"  ;
    if (arc_index == 1710) return "W"  ;
    if (arc_index == 1711) return "W"  ;
    if (arc_index == 1712) return "W"  ;
    if (arc_index == 1713) return "W"  ;
    if (arc_index == 1714) return "E"  ;
    if (arc_index == 1715) return "W"  ;
    if (arc_index == 1727) return "H"  ;
    if (arc_index == 1761) return "H"  ;
    if (arc_index == 1762) return "W"  ;
    if (arc_index == 1767) return "W"  ;
    if (arc_index == 1771) return "W"  ;
    if (arc_index == 1772) return "H"  ;
    if (arc_index == 1838) return "E"  ;
    if (arc_index == 1946) return "E"  ;
    if (arc_index == 1971) return "H"  ;
    if (arc_index == 2037) return "E"  ;
    if (arc_index == 2094) return "W"  ;
    if (arc_index == 2102) return "W"  ;
    if (arc_index == 2110) return "W"  ;
    if (arc_index == 2148) return "H"  ;
    if (arc_index == 2232) return "H"  ;
    if (arc_index == 2265) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2335) return "W"  ;
    if (arc_index == 2341) return "H"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2457) return "H"  ;
    if (arc_index == 2530) return "W"  ;
    if (arc_index == 2544) return "E"  ;
    if (arc_index == 2546) return "H"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2558) return "E"  ;
    if (arc_index == 2560) return "H"  ;
    if (arc_index == 2563) return "H"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2691) return "H"  ;
    if (arc_index == 2732) return "E"  ;
    if (arc_index == 2737) return "E"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2776) return "E"  ;
    if (arc_index == 2777) return "E"  ;
    if (arc_index == 2779) return "E"  ;
    if (arc_index == 2786) return "E"  ;
    if (arc_index == 2790) return "E"  ;
    if (arc_index == 2791) return "E"  ;
    if (arc_index == 2829) return "W"  ;
    if (arc_index == 2844) return "H"  ;
    if (arc_index == 2853) return "E"  ;
    if (arc_index == 2858) return "E"  ;
    if (arc_index == 2916) return "W"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 2)) begin 
    if (arc_index == 41) return "W"  ;
    if (arc_index == 49) return "W"  ;
    if (arc_index == 80) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 115) return "W"  ;
    if (arc_index == 136) return "W"  ;
    if (arc_index == 202) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 244) return "W"  ;
    if (arc_index == 247) return "W"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 443) return "W"  ;
    if (arc_index == 550) return "W"  ;
    if (arc_index == 571) return "W"  ;
    if (arc_index == 577) return "E"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 587) return "E"  ;
    if (arc_index == 589) return "H"  ;
    if (arc_index == 654) return "W"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 744) return "H"  ;
    if (arc_index == 751) return "H"  ;
    if (arc_index == 753) return "W"  ;
    if (arc_index == 761) return "W"  ;
    if (arc_index == 770) return "W"  ;
    if (arc_index == 779) return "W"  ;
    if (arc_index == 787) return "W"  ;
    if (arc_index == 789) return "W"  ;
    if (arc_index == 799) return "W"  ;
    if (arc_index == 803) return "W"  ;
    if (arc_index == 816) return "W"  ;
    if (arc_index == 840) return "W"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 877) return "H"  ;
    if (arc_index == 880) return "H"  ;
    if (arc_index == 882) return "E"  ;
    if (arc_index == 884) return "E"  ;
    if (arc_index == 885) return "H"  ;
    if (arc_index == 886) return "H"  ;
    if (arc_index == 888) return "H"  ;
    if (arc_index == 890) return "E"  ;
    if (arc_index == 894) return "W"  ;
    if (arc_index == 895) return "E"  ;
    if (arc_index == 896) return "E"  ;
    if (arc_index == 898) return "E"  ;
    if (arc_index == 900) return "E"  ;
    if (arc_index == 907) return "E"  ;
    if (arc_index == 913) return "E"  ;
    if (arc_index == 931) return "W"  ;
    if (arc_index == 949) return "E"  ;
    if (arc_index == 951) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 958) return "E"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 961) return "E"  ;
    if (arc_index == 967) return "E"  ;
    if (arc_index == 972) return "H"  ;
    if (arc_index == 994) return "H"  ;
    if (arc_index == 1056) return "W"  ;
    if (arc_index == 1078) return "E"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1082) return "E"  ;
    if (arc_index == 1083) return "E"  ;
    if (arc_index == 1085) return "E"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1088) return "E"  ;
    if (arc_index == 1089) return "E"  ;
    if (arc_index == 1091) return "E"  ;
    if (arc_index == 1092) return "E"  ;
    if (arc_index == 1093) return "E"  ;
    if (arc_index == 1094) return "E"  ;
    if (arc_index == 1098) return "H"  ;
    if (arc_index == 1111) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1193) return "E"  ;
    if (arc_index == 1202) return "E"  ;
    if (arc_index == 1209) return "H"  ;
    if (arc_index == 1224) return "H"  ;
    if (arc_index == 1231) return "H"  ;
    if (arc_index == 1279) return "H"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1400) return "W"  ;
    if (arc_index == 1454) return "H"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1484) return "W"  ;
    if (arc_index == 1527) return "W"  ;
    if (arc_index == 1533) return "W"  ;
    if (arc_index == 1616) return "W"  ;
    if (arc_index == 1636) return "W"  ;
    if (arc_index == 1643) return "W"  ;
    if (arc_index == 1647) return "E"  ;
    if (arc_index == 1651) return "H"  ;
    if (arc_index == 1673) return "H"  ;
    if (arc_index == 1694) return "H"  ;
    if (arc_index == 1706) return "H"  ;
    if (arc_index == 1709) return "W"  ;
    if (arc_index == 1716) return "W"  ;
    if (arc_index == 1717) return "E"  ;
    if (arc_index == 1718) return "E"  ;
    if (arc_index == 1719) return "E"  ;
    if (arc_index == 1720) return "E"  ;
    if (arc_index == 1721) return "E"  ;
    if (arc_index == 1722) return "W"  ;
    if (arc_index == 1723) return "W"  ;
    if (arc_index == 1724) return "E"  ;
    if (arc_index == 1725) return "W"  ;
    if (arc_index == 1726) return "W"  ;
    if (arc_index == 1727) return "E"  ;
    if (arc_index == 1728) return "E"  ;
    if (arc_index == 1729) return "E"  ;
    if (arc_index == 1730) return "E"  ;
    if (arc_index == 1731) return "E"  ;
    if (arc_index == 1732) return "E"  ;
    if (arc_index == 1733) return "W"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1735) return "E"  ;
    if (arc_index == 1736) return "E"  ;
    if (arc_index == 1737) return "E"  ;
    if (arc_index == 1740) return "E"  ;
    if (arc_index == 1743) return "E"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1749) return "H"  ;
    if (arc_index == 1752) return "H"  ;
    if (arc_index == 1753) return "E"  ;
    if (arc_index == 1754) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1768) return "E"  ;
    if (arc_index == 1794) return "H"  ;
    if (arc_index == 1798) return "W"  ;
    if (arc_index == 1808) return "W"  ;
    if (arc_index == 1812) return "W"  ;
    if (arc_index == 1841) return "W"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1897) return "W"  ;
    if (arc_index == 1915) return "E"  ;
    if (arc_index == 1919) return "E"  ;
    if (arc_index == 1920) return "E"  ;
    if (arc_index == 1933) return "E"  ;
    if (arc_index == 1934) return "W"  ;
    if (arc_index == 1963) return "W"  ;
    if (arc_index == 1993) return "H"  ;
    if (arc_index == 2002) return "E"  ;
    if (arc_index == 2015) return "E"  ;
    if (arc_index == 2038) return "W"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2170) return "H"  ;
    if (arc_index == 2254) return "H"  ;
    if (arc_index == 2276) return "H"  ;
    if (arc_index == 2305) return "W"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2363) return "H"  ;
    if (arc_index == 2474) return "W"  ;
    if (arc_index == 2479) return "H"  ;
    if (arc_index == 2480) return "H"  ;
    if (arc_index == 2557) return "H"  ;
    if (arc_index == 2568) return "H"  ;
    if (arc_index == 2576) return "E"  ;
    if (arc_index == 2582) return "H"  ;
    if (arc_index == 2590) return "H"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2679) return "E"  ;
    if (arc_index == 2713) return "H"  ;
    if (arc_index == 2760) return "H"  ;
    if (arc_index == 2761) return "W"  ;
    if (arc_index == 2765) return "W"  ;
    if (arc_index == 2780) return "W"  ;
    if (arc_index == 2788) return "W"  ;
    if (arc_index == 2792) return "W"  ;
    if (arc_index == 2800) return "E"  ;
    if (arc_index == 2803) return "E"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2809) return "E"  ;
    if (arc_index == 2834) return "E"  ;
    if (arc_index == 2861) return "E"  ;
    if (arc_index == 2866) return "H"  ;
    if (arc_index == 2875) return "H"  ;
    if (arc_index == 2900) return "W"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 2)) begin 
    if (arc_index == 12) return "W"  ;
    if (arc_index == 80) return "W"  ;
    if (arc_index == 152) return "W"  ;
    if (arc_index == 211) return "W"  ;
    if (arc_index == 256) return "W"  ;
    if (arc_index == 340) return "W"  ;
    if (arc_index == 472) return "W"  ;
    if (arc_index == 486) return "E"  ;
    if (arc_index == 493) return "E"  ;
    if (arc_index == 508) return "E"  ;
    if (arc_index == 611) return "H"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 766) return "H"  ;
    if (arc_index == 770) return "H"  ;
    if (arc_index == 774) return "H"  ;
    if (arc_index == 779) return "H"  ;
    if (arc_index == 783) return "H"  ;
    if (arc_index == 787) return "H"  ;
    if (arc_index == 789) return "H"  ;
    if (arc_index == 803) return "H"  ;
    if (arc_index == 848) return "H"  ;
    if (arc_index == 889) return "E"  ;
    if (arc_index == 897) return "E"  ;
    if (arc_index == 899) return "H"  ;
    if (arc_index == 907) return "H"  ;
    if (arc_index == 950) return "E"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 994) return "H"  ;
    if (arc_index == 1120) return "H"  ;
    if (arc_index == 1202) return "E"  ;
    if (arc_index == 1224) return "E"  ;
    if (arc_index == 1231) return "H"  ;
    if (arc_index == 1301) return "H"  ;
    if (arc_index == 1418) return "H"  ;
    if (arc_index == 1424) return "H"  ;
    if (arc_index == 1454) return "H"  ;
    if (arc_index == 1476) return "H"  ;
    if (arc_index == 1533) return "H"  ;
    if (arc_index == 1600) return "E"  ;
    if (arc_index == 1622) return "E"  ;
    if (arc_index == 1636) return "E"  ;
    if (arc_index == 1673) return "H"  ;
    if (arc_index == 1706) return "H"  ;
    if (arc_index == 1709) return "H"  ;
    if (arc_index == 1716) return "H"  ;
    if (arc_index == 1721) return "H"  ;
    if (arc_index == 1738) return "E"  ;
    if (arc_index == 1739) return "E"  ;
    if (arc_index == 1740) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1742) return "E"  ;
    if (arc_index == 1743) return "E"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1745) return "E"  ;
    if (arc_index == 1746) return "E"  ;
    if (arc_index == 1747) return "E"  ;
    if (arc_index == 1748) return "E"  ;
    if (arc_index == 1749) return "E"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1751) return "E"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1753) return "E"  ;
    if (arc_index == 1754) return "E"  ;
    if (arc_index == 1755) return "E"  ;
    if (arc_index == 1756) return "W"  ;
    if (arc_index == 1757) return "E"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1771) return "H"  ;
    if (arc_index == 1816) return "H"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1920) return "W"  ;
    if (arc_index == 1984) return "W"  ;
    if (arc_index == 2015) return "H"  ;
    if (arc_index == 2029) return "W"  ;
    if (arc_index == 2030) return "W"  ;
    if (arc_index == 2192) return "H"  ;
    if (arc_index == 2232) return "H"  ;
    if (arc_index == 2276) return "H"  ;
    if (arc_index == 2291) return "W"  ;
    if (arc_index == 2305) return "W"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2385) return "H"  ;
    if (arc_index == 2466) return "W"  ;
    if (arc_index == 2501) return "H"  ;
    if (arc_index == 2562) return "E"  ;
    if (arc_index == 2564) return "E"  ;
    if (arc_index == 2568) return "E"  ;
    if (arc_index == 2590) return "H"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2604) return "H"  ;
    if (arc_index == 2671) return "E"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2728) return "E"  ;
    if (arc_index == 2731) return "E"  ;
    if (arc_index == 2732) return "E"  ;
    if (arc_index == 2735) return "H"  ;
    if (arc_index == 2736) return "E"  ;
    if (arc_index == 2737) return "E"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2742) return "E"  ;
    if (arc_index == 2744) return "E"  ;
    if (arc_index == 2749) return "E"  ;
    if (arc_index == 2838) return "W"  ;
    if (arc_index == 2851) return "W"  ;
    if (arc_index == 2861) return "W"  ;
    if (arc_index == 2862) return "W"  ;
    if (arc_index == 2864) return "E"  ;
    if (arc_index == 2865) return "E"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2871) return "E"  ;
    if (arc_index == 2873) return "E"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2876) return "E"  ;
    if (arc_index == 2888) return "H"  ;
    if (arc_index == 2893) return "W"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 9)) begin 
    if (arc_index == 314) return "W"  ;
    if (arc_index == 551) return "E"  ;
    if (arc_index == 558) return "E"  ;
    if (arc_index == 563) return "E"  ;
    if (arc_index == 628) return "W"  ;
    if (arc_index == 633) return "H"  ;
    if (arc_index == 788) return "H"  ;
    if (arc_index == 921) return "H"  ;
    if (arc_index == 929) return "H"  ;
    if (arc_index == 1016) return "H"  ;
    if (arc_index == 1142) return "H"  ;
    if (arc_index == 1253) return "H"  ;
    if (arc_index == 1323) return "H"  ;
    if (arc_index == 1343) return "W"  ;
    if (arc_index == 1346) return "W"  ;
    if (arc_index == 1498) return "H"  ;
    if (arc_index == 1547) return "W"  ;
    if (arc_index == 1695) return "H"  ;
    if (arc_index == 1738) return "H"  ;
    if (arc_index == 1760) return "W"  ;
    if (arc_index == 1761) return "W"  ;
    if (arc_index == 1762) return "W"  ;
    if (arc_index == 1763) return "W"  ;
    if (arc_index == 1764) return "W"  ;
    if (arc_index == 1765) return "W"  ;
    if (arc_index == 1766) return "E"  ;
    if (arc_index == 1767) return "W"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1769) return "W"  ;
    if (arc_index == 1770) return "W"  ;
    if (arc_index == 1771) return "W"  ;
    if (arc_index == 1772) return "W"  ;
    if (arc_index == 1773) return "W"  ;
    if (arc_index == 1774) return "W"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1777) return "E"  ;
    if (arc_index == 1778) return "W"  ;
    if (arc_index == 1779) return "E"  ;
    if (arc_index == 1780) return "E"  ;
    if (arc_index == 1781) return "W"  ;
    if (arc_index == 1793) return "H"  ;
    if (arc_index == 1838) return "H"  ;
    if (arc_index == 2037) return "H"  ;
    if (arc_index == 2101) return "E"  ;
    if (arc_index == 2105) return "E"  ;
    if (arc_index == 2107) return "E"  ;
    if (arc_index == 2111) return "E"  ;
    if (arc_index == 2214) return "H"  ;
    if (arc_index == 2298) return "H"  ;
    if (arc_index == 2349) return "W"  ;
    if (arc_index == 2407) return "H"  ;
    if (arc_index == 2523) return "H"  ;
    if (arc_index == 2612) return "H"  ;
    if (arc_index == 2626) return "H"  ;
    if (arc_index == 2628) return "W"  ;
    if (arc_index == 2757) return "H"  ;
    if (arc_index == 2910) return "H"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 6)) begin 
    if (arc_index == 4) return "H"  ;
    if (arc_index == 5) return "H"  ;
    if (arc_index == 6) return "H"  ;
    if (arc_index == 9) return "H"  ;
    if (arc_index == 12) return "W"  ;
    if (arc_index == 14) return "W"  ;
    if (arc_index == 16) return "E"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 113) return "E"  ;
    if (arc_index == 125) return "E"  ;
    if (arc_index == 202) return "W"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 212) return "W"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 261) return "W"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 278) return "W"  ;
    if (arc_index == 301) return "W"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 340) return "W"  ;
    if (arc_index == 399) return "W"  ;
    if (arc_index == 403) return "W"  ;
    if (arc_index == 426) return "W"  ;
    if (arc_index == 436) return "W"  ;
    if (arc_index == 442) return "W"  ;
    if (arc_index == 475) return "W"  ;
    if (arc_index == 480) return "W"  ;
    if (arc_index == 485) return "W"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 512) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 547) return "E"  ;
    if (arc_index == 557) return "W"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 613) return "W"  ;
    if (arc_index == 634) return "W"  ;
    if (arc_index == 642) return "W"  ;
    if (arc_index == 655) return "H"  ;
    if (arc_index == 690) return "W"  ;
    if (arc_index == 691) return "W"  ;
    if (arc_index == 693) return "W"  ;
    if (arc_index == 710) return "W"  ;
    if (arc_index == 719) return "W"  ;
    if (arc_index == 756) return "E"  ;
    if (arc_index == 763) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 810) return "H"  ;
    if (arc_index == 815) return "W"  ;
    if (arc_index == 816) return "W"  ;
    if (arc_index == 819) return "W"  ;
    if (arc_index == 821) return "W"  ;
    if (arc_index == 822) return "W"  ;
    if (arc_index == 826) return "W"  ;
    if (arc_index == 836) return "W"  ;
    if (arc_index == 837) return "W"  ;
    if (arc_index == 838) return "W"  ;
    if (arc_index == 839) return "W"  ;
    if (arc_index == 850) return "W"  ;
    if (arc_index == 851) return "W"  ;
    if (arc_index == 852) return "W"  ;
    if (arc_index == 857) return "W"  ;
    if (arc_index == 863) return "W"  ;
    if (arc_index == 869) return "W"  ;
    if (arc_index == 883) return "W"  ;
    if (arc_index == 887) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 943) return "H"  ;
    if (arc_index == 945) return "H"  ;
    if (arc_index == 951) return "H"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 967) return "E"  ;
    if (arc_index == 971) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1038) return "H"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1062) return "W"  ;
    if (arc_index == 1076) return "W"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1088) return "E"  ;
    if (arc_index == 1089) return "E"  ;
    if (arc_index == 1091) return "E"  ;
    if (arc_index == 1108) return "E"  ;
    if (arc_index == 1113) return "E"  ;
    if (arc_index == 1120) return "E"  ;
    if (arc_index == 1124) return "E"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1164) return "H"  ;
    if (arc_index == 1174) return "H"  ;
    if (arc_index == 1187) return "W"  ;
    if (arc_index == 1190) return "W"  ;
    if (arc_index == 1220) return "W"  ;
    if (arc_index == 1236) return "W"  ;
    if (arc_index == 1257) return "W"  ;
    if (arc_index == 1275) return "H"  ;
    if (arc_index == 1286) return "H"  ;
    if (arc_index == 1290) return "H"  ;
    if (arc_index == 1334) return "H"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1345) return "H"  ;
    if (arc_index == 1349) return "H"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1359) return "W"  ;
    if (arc_index == 1362) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1394) return "W"  ;
    if (arc_index == 1396) return "W"  ;
    if (arc_index == 1398) return "W"  ;
    if (arc_index == 1401) return "W"  ;
    if (arc_index == 1405) return "W"  ;
    if (arc_index == 1410) return "E"  ;
    if (arc_index == 1413) return "E"  ;
    if (arc_index == 1415) return "E"  ;
    if (arc_index == 1421) return "E"  ;
    if (arc_index == 1422) return "E"  ;
    if (arc_index == 1423) return "E"  ;
    if (arc_index == 1449) return "E"  ;
    if (arc_index == 1452) return "E"  ;
    if (arc_index == 1455) return "W"  ;
    if (arc_index == 1456) return "W"  ;
    if (arc_index == 1461) return "E"  ;
    if (arc_index == 1462) return "E"  ;
    if (arc_index == 1470) return "E"  ;
    if (arc_index == 1471) return "E"  ;
    if (arc_index == 1477) return "W"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1483) return "W"  ;
    if (arc_index == 1484) return "W"  ;
    if (arc_index == 1485) return "W"  ;
    if (arc_index == 1492) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1520) return "H"  ;
    if (arc_index == 1530) return "H"  ;
    if (arc_index == 1534) return "H"  ;
    if (arc_index == 1543) return "H"  ;
    if (arc_index == 1580) return "H"  ;
    if (arc_index == 1624) return "H"  ;
    if (arc_index == 1666) return "E"  ;
    if (arc_index == 1703) return "E"  ;
    if (arc_index == 1704) return "E"  ;
    if (arc_index == 1717) return "H"  ;
    if (arc_index == 1736) return "H"  ;
    if (arc_index == 1744) return "H"  ;
    if (arc_index == 1751) return "E"  ;
    if (arc_index == 1760) return "H"  ;
    if (arc_index == 1773) return "H"  ;
    if (arc_index == 1776) return "H"  ;
    if (arc_index == 1778) return "W"  ;
    if (arc_index == 1782) return "W"  ;
    if (arc_index == 1783) return "W"  ;
    if (arc_index == 1784) return "W"  ;
    if (arc_index == 1785) return "W"  ;
    if (arc_index == 1786) return "W"  ;
    if (arc_index == 1787) return "W"  ;
    if (arc_index == 1788) return "W"  ;
    if (arc_index == 1789) return "W"  ;
    if (arc_index == 1790) return "W"  ;
    if (arc_index == 1791) return "E"  ;
    if (arc_index == 1792) return "E"  ;
    if (arc_index == 1793) return "E"  ;
    if (arc_index == 1794) return "W"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1796) return "E"  ;
    if (arc_index == 1797) return "E"  ;
    if (arc_index == 1798) return "W"  ;
    if (arc_index == 1799) return "W"  ;
    if (arc_index == 1800) return "W"  ;
    if (arc_index == 1801) return "W"  ;
    if (arc_index == 1802) return "W"  ;
    if (arc_index == 1803) return "W"  ;
    if (arc_index == 1808) return "W"  ;
    if (arc_index == 1815) return "H"  ;
    if (arc_index == 1832) return "E"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1837) return "E"  ;
    if (arc_index == 1844) return "E"  ;
    if (arc_index == 1847) return "E"  ;
    if (arc_index == 1852) return "E"  ;
    if (arc_index == 1860) return "H"  ;
    if (arc_index == 1862) return "H"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1906) return "W"  ;
    if (arc_index == 1928) return "E"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1958) return "W"  ;
    if (arc_index == 1959) return "W"  ;
    if (arc_index == 1963) return "W"  ;
    if (arc_index == 1971) return "W"  ;
    if (arc_index == 1979) return "W"  ;
    if (arc_index == 1985) return "E"  ;
    if (arc_index == 1989) return "E"  ;
    if (arc_index == 1991) return "E"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 1996) return "E"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2055) return "E"  ;
    if (arc_index == 2059) return "H"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2091) return "E"  ;
    if (arc_index == 2097) return "E"  ;
    if (arc_index == 2103) return "W"  ;
    if (arc_index == 2123) return "E"  ;
    if (arc_index == 2152) return "E"  ;
    if (arc_index == 2171) return "E"  ;
    if (arc_index == 2236) return "H"  ;
    if (arc_index == 2252) return "H"  ;
    if (arc_index == 2260) return "H"  ;
    if (arc_index == 2262) return "H"  ;
    if (arc_index == 2265) return "H"  ;
    if (arc_index == 2268) return "H"  ;
    if (arc_index == 2274) return "H"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2302) return "W"  ;
    if (arc_index == 2318) return "W"  ;
    if (arc_index == 2320) return "H"  ;
    if (arc_index == 2346) return "H"  ;
    if (arc_index == 2364) return "W"  ;
    if (arc_index == 2429) return "H"  ;
    if (arc_index == 2449) return "H"  ;
    if (arc_index == 2468) return "H"  ;
    if (arc_index == 2470) return "E"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2490) return "E"  ;
    if (arc_index == 2492) return "E"  ;
    if (arc_index == 2496) return "E"  ;
    if (arc_index == 2503) return "E"  ;
    if (arc_index == 2504) return "E"  ;
    if (arc_index == 2506) return "E"  ;
    if (arc_index == 2543) return "E"  ;
    if (arc_index == 2545) return "H"  ;
    if (arc_index == 2548) return "H"  ;
    if (arc_index == 2554) return "E"  ;
    if (arc_index == 2567) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2611) return "W"  ;
    if (arc_index == 2634) return "H"  ;
    if (arc_index == 2648) return "H"  ;
    if (arc_index == 2687) return "H"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2751) return "E"  ;
    if (arc_index == 2753) return "E"  ;
    if (arc_index == 2768) return "E"  ;
    if (arc_index == 2769) return "E"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2779) return "H"  ;
    if (arc_index == 2782) return "H"  ;
    if (arc_index == 2794) return "E"  ;
    if (arc_index == 2810) return "E"  ;
    if (arc_index == 2823) return "W"  ;
    if (arc_index == 2827) return "W"  ;
    if (arc_index == 2828) return "W"  ;
    if (arc_index == 2834) return "W"  ;
    if (arc_index == 2835) return "W"  ;
    if (arc_index == 2849) return "E"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2855) return "E"  ;
    if (arc_index == 2882) return "E"  ;
    if (arc_index == 2894) return "E"  ;
    if (arc_index == 2901) return "E"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2918) return "W"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 7)) begin 
    if (arc_index == 28) return "H"  ;
    if (arc_index == 30) return "H"  ;
    if (arc_index == 43) return "H"  ;
    if (arc_index == 92) return "H"  ;
    if (arc_index == 95) return "H"  ;
    if (arc_index == 133) return "H"  ;
    if (arc_index == 158) return "W"  ;
    if (arc_index == 159) return "W"  ;
    if (arc_index == 160) return "W"  ;
    if (arc_index == 176) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 198) return "W"  ;
    if (arc_index == 201) return "W"  ;
    if (arc_index == 206) return "W"  ;
    if (arc_index == 209) return "W"  ;
    if (arc_index == 210) return "W"  ;
    if (arc_index == 217) return "W"  ;
    if (arc_index == 219) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 276) return "W"  ;
    if (arc_index == 278) return "W"  ;
    if (arc_index == 281) return "W"  ;
    if (arc_index == 288) return "W"  ;
    if (arc_index == 308) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 312) return "W"  ;
    if (arc_index == 315) return "W"  ;
    if (arc_index == 327) return "W"  ;
    if (arc_index == 344) return "W"  ;
    if (arc_index == 347) return "E"  ;
    if (arc_index == 354) return "E"  ;
    if (arc_index == 359) return "E"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 428) return "E"  ;
    if (arc_index == 433) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 537) return "E"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 554) return "W"  ;
    if (arc_index == 561) return "W"  ;
    if (arc_index == 564) return "W"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 649) return "W"  ;
    if (arc_index == 652) return "W"  ;
    if (arc_index == 653) return "W"  ;
    if (arc_index == 677) return "H"  ;
    if (arc_index == 686) return "W"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 721) return "W"  ;
    if (arc_index == 736) return "W"  ;
    if (arc_index == 742) return "W"  ;
    if (arc_index == 758) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 831) return "E"  ;
    if (arc_index == 832) return "H"  ;
    if (arc_index == 841) return "E"  ;
    if (arc_index == 857) return "E"  ;
    if (arc_index == 882) return "E"  ;
    if (arc_index == 883) return "E"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 965) return "H"  ;
    if (arc_index == 973) return "H"  ;
    if (arc_index == 981) return "H"  ;
    if (arc_index == 1050) return "H"  ;
    if (arc_index == 1052) return "H"  ;
    if (arc_index == 1060) return "H"  ;
    if (arc_index == 1064) return "H"  ;
    if (arc_index == 1070) return "H"  ;
    if (arc_index == 1076) return "H"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1103) return "E"  ;
    if (arc_index == 1118) return "E"  ;
    if (arc_index == 1147) return "E"  ;
    if (arc_index == 1149) return "W"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1161) return "W"  ;
    if (arc_index == 1164) return "W"  ;
    if (arc_index == 1186) return "H"  ;
    if (arc_index == 1195) return "H"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1257) return "E"  ;
    if (arc_index == 1286) return "W"  ;
    if (arc_index == 1297) return "H"  ;
    if (arc_index == 1313) return "H"  ;
    if (arc_index == 1321) return "H"  ;
    if (arc_index == 1334) return "W"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1341) return "W"  ;
    if (arc_index == 1344) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1367) return "H"  ;
    if (arc_index == 1374) return "H"  ;
    if (arc_index == 1379) return "H"  ;
    if (arc_index == 1394) return "E"  ;
    if (arc_index == 1398) return "E"  ;
    if (arc_index == 1399) return "E"  ;
    if (arc_index == 1427) return "E"  ;
    if (arc_index == 1460) return "E"  ;
    if (arc_index == 1494) return "E"  ;
    if (arc_index == 1515) return "E"  ;
    if (arc_index == 1541) return "W"  ;
    if (arc_index == 1542) return "H"  ;
    if (arc_index == 1543) return "W"  ;
    if (arc_index == 1554) return "W"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1610) return "E"  ;
    if (arc_index == 1613) return "E"  ;
    if (arc_index == 1619) return "E"  ;
    if (arc_index == 1653) return "E"  ;
    if (arc_index == 1654) return "E"  ;
    if (arc_index == 1689) return "E"  ;
    if (arc_index == 1736) return "E"  ;
    if (arc_index == 1739) return "H"  ;
    if (arc_index == 1764) return "H"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1782) return "H"  ;
    if (arc_index == 1787) return "E"  ;
    if (arc_index == 1792) return "E"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1803) return "E"  ;
    if (arc_index == 1804) return "W"  ;
    if (arc_index == 1805) return "E"  ;
    if (arc_index == 1806) return "E"  ;
    if (arc_index == 1807) return "E"  ;
    if (arc_index == 1808) return "W"  ;
    if (arc_index == 1809) return "E"  ;
    if (arc_index == 1810) return "E"  ;
    if (arc_index == 1811) return "E"  ;
    if (arc_index == 1812) return "W"  ;
    if (arc_index == 1813) return "W"  ;
    if (arc_index == 1814) return "W"  ;
    if (arc_index == 1815) return "W"  ;
    if (arc_index == 1816) return "W"  ;
    if (arc_index == 1817) return "E"  ;
    if (arc_index == 1818) return "E"  ;
    if (arc_index == 1819) return "E"  ;
    if (arc_index == 1820) return "E"  ;
    if (arc_index == 1821) return "E"  ;
    if (arc_index == 1822) return "W"  ;
    if (arc_index == 1823) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1825) return "E"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1837) return "H"  ;
    if (arc_index == 1847) return "E"  ;
    if (arc_index == 1851) return "E"  ;
    if (arc_index == 1858) return "E"  ;
    if (arc_index == 1867) return "E"  ;
    if (arc_index == 1869) return "E"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1882) return "H"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1917) return "E"  ;
    if (arc_index == 1958) return "E"  ;
    if (arc_index == 1959) return "E"  ;
    if (arc_index == 1963) return "E"  ;
    if (arc_index == 1971) return "E"  ;
    if (arc_index == 1977) return "E"  ;
    if (arc_index == 1978) return "E"  ;
    if (arc_index == 1991) return "E"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2081) return "H"  ;
    if (arc_index == 2090) return "W"  ;
    if (arc_index == 2095) return "W"  ;
    if (arc_index == 2121) return "E"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2215) return "E"  ;
    if (arc_index == 2237) return "E"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2258) return "H"  ;
    if (arc_index == 2266) return "H"  ;
    if (arc_index == 2268) return "W"  ;
    if (arc_index == 2285) return "W"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2288) return "W"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2294) return "E"  ;
    if (arc_index == 2296) return "E"  ;
    if (arc_index == 2299) return "E"  ;
    if (arc_index == 2303) return "E"  ;
    if (arc_index == 2306) return "E"  ;
    if (arc_index == 2307) return "E"  ;
    if (arc_index == 2308) return "W"  ;
    if (arc_index == 2313) return "W"  ;
    if (arc_index == 2318) return "W"  ;
    if (arc_index == 2321) return "W"  ;
    if (arc_index == 2342) return "H"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2363) return "W"  ;
    if (arc_index == 2366) return "W"  ;
    if (arc_index == 2368) return "W"  ;
    if (arc_index == 2369) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2375) return "W"  ;
    if (arc_index == 2386) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2413) return "W"  ;
    if (arc_index == 2424) return "W"  ;
    if (arc_index == 2432) return "E"  ;
    if (arc_index == 2451) return "H"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2470) return "E"  ;
    if (arc_index == 2476) return "E"  ;
    if (arc_index == 2482) return "E"  ;
    if (arc_index == 2496) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2538) return "E"  ;
    if (arc_index == 2548) return "E"  ;
    if (arc_index == 2567) return "H"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2605) return "W"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2620) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2627) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2656) return "H"  ;
    if (arc_index == 2670) return "H"  ;
    if (arc_index == 2703) return "H"  ;
    if (arc_index == 2714) return "W"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2801) return "H"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2810) return "E"  ;
    if (arc_index == 2817) return "W"  ;
    if (arc_index == 2819) return "W"  ;
    if (arc_index == 2820) return "W"  ;
    if (arc_index == 2821) return "W"  ;
    if (arc_index == 2822) return "E"  ;
    if (arc_index == 2824) return "E"  ;
    if (arc_index == 2825) return "E"  ;
    if (arc_index == 2831) return "E"  ;
    if (arc_index == 2837) return "E"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2855) return "E"  ;
    if (arc_index == 2892) return "E"  ;
    if (arc_index == 2912) return "E"  ;
    if (arc_index == 2915) return "E"  ;
    if (arc_index == 2919) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 3)) begin 
    if (arc_index == 26) return "W"  ;
    if (arc_index == 41) return "W"  ;
    if (arc_index == 49) return "W"  ;
    if (arc_index == 50) return "H"  ;
    if (arc_index == 76) return "H"  ;
    if (arc_index == 152) return "H"  ;
    if (arc_index == 200) return "H"  ;
    if (arc_index == 202) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 384) return "W"  ;
    if (arc_index == 390) return "W"  ;
    if (arc_index == 404) return "W"  ;
    if (arc_index == 470) return "E"  ;
    if (arc_index == 471) return "E"  ;
    if (arc_index == 472) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 570) return "E"  ;
    if (arc_index == 571) return "W"  ;
    if (arc_index == 574) return "E"  ;
    if (arc_index == 577) return "E"  ;
    if (arc_index == 587) return "E"  ;
    if (arc_index == 664) return "E"  ;
    if (arc_index == 675) return "E"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 699) return "H"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 750) return "W"  ;
    if (arc_index == 755) return "W"  ;
    if (arc_index == 761) return "W"  ;
    if (arc_index == 785) return "W"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 816) return "W"  ;
    if (arc_index == 854) return "H"  ;
    if (arc_index == 882) return "E"  ;
    if (arc_index == 890) return "E"  ;
    if (arc_index == 895) return "E"  ;
    if (arc_index == 909) return "E"  ;
    if (arc_index == 914) return "E"  ;
    if (arc_index == 949) return "E"  ;
    if (arc_index == 951) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 961) return "E"  ;
    if (arc_index == 967) return "E"  ;
    if (arc_index == 972) return "W"  ;
    if (arc_index == 987) return "H"  ;
    if (arc_index == 995) return "H"  ;
    if (arc_index == 1078) return "E"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1082) return "H"  ;
    if (arc_index == 1085) return "H"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1088) return "E"  ;
    if (arc_index == 1089) return "E"  ;
    if (arc_index == 1091) return "E"  ;
    if (arc_index == 1092) return "E"  ;
    if (arc_index == 1093) return "E"  ;
    if (arc_index == 1094) return "E"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1193) return "W"  ;
    if (arc_index == 1208) return "H"  ;
    if (arc_index == 1279) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1319) return "H"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1389) return "H"  ;
    if (arc_index == 1407) return "H"  ;
    if (arc_index == 1465) return "H"  ;
    if (arc_index == 1477) return "H"  ;
    if (arc_index == 1478) return "H"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1484) return "W"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1564) return "H"  ;
    if (arc_index == 1587) return "H"  ;
    if (arc_index == 1599) return "H"  ;
    if (arc_index == 1622) return "H"  ;
    if (arc_index == 1629) return "H"  ;
    if (arc_index == 1633) return "H"  ;
    if (arc_index == 1647) return "E"  ;
    if (arc_index == 1651) return "W"  ;
    if (arc_index == 1667) return "W"  ;
    if (arc_index == 1694) return "W"  ;
    if (arc_index == 1712) return "W"  ;
    if (arc_index == 1715) return "W"  ;
    if (arc_index == 1717) return "E"  ;
    if (arc_index == 1724) return "E"  ;
    if (arc_index == 1727) return "E"  ;
    if (arc_index == 1728) return "E"  ;
    if (arc_index == 1730) return "E"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1736) return "E"  ;
    if (arc_index == 1737) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1753) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1761) return "H"  ;
    if (arc_index == 1794) return "W"  ;
    if (arc_index == 1798) return "W"  ;
    if (arc_index == 1804) return "H"  ;
    if (arc_index == 1808) return "W"  ;
    if (arc_index == 1812) return "W"  ;
    if (arc_index == 1822) return "W"  ;
    if (arc_index == 1826) return "E"  ;
    if (arc_index == 1827) return "E"  ;
    if (arc_index == 1828) return "E"  ;
    if (arc_index == 1829) return "E"  ;
    if (arc_index == 1830) return "E"  ;
    if (arc_index == 1831) return "E"  ;
    if (arc_index == 1832) return "E"  ;
    if (arc_index == 1833) return "E"  ;
    if (arc_index == 1834) return "E"  ;
    if (arc_index == 1835) return "E"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1837) return "E"  ;
    if (arc_index == 1838) return "E"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1840) return "E"  ;
    if (arc_index == 1841) return "W"  ;
    if (arc_index == 1842) return "W"  ;
    if (arc_index == 1843) return "W"  ;
    if (arc_index == 1844) return "E"  ;
    if (arc_index == 1845) return "E"  ;
    if (arc_index == 1846) return "E"  ;
    if (arc_index == 1847) return "E"  ;
    if (arc_index == 1859) return "H"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1904) return "H"  ;
    if (arc_index == 1915) return "E"  ;
    if (arc_index == 1919) return "E"  ;
    if (arc_index == 1933) return "E"  ;
    if (arc_index == 1941) return "E"  ;
    if (arc_index == 1963) return "W"  ;
    if (arc_index == 1987) return "W"  ;
    if (arc_index == 1992) return "W"  ;
    if (arc_index == 2001) return "W"  ;
    if (arc_index == 2002) return "W"  ;
    if (arc_index == 2007) return "W"  ;
    if (arc_index == 2024) return "W"  ;
    if (arc_index == 2032) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2035) return "E"  ;
    if (arc_index == 2036) return "E"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2040) return "E"  ;
    if (arc_index == 2042) return "E"  ;
    if (arc_index == 2043) return "E"  ;
    if (arc_index == 2050) return "E"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2103) return "H"  ;
    if (arc_index == 2170) return "W"  ;
    if (arc_index == 2171) return "E"  ;
    if (arc_index == 2202) return "E"  ;
    if (arc_index == 2254) return "W"  ;
    if (arc_index == 2276) return "W"  ;
    if (arc_index == 2280) return "H"  ;
    if (arc_index == 2297) return "H"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2363) return "W"  ;
    if (arc_index == 2364) return "H"  ;
    if (arc_index == 2399) return "H"  ;
    if (arc_index == 2434) return "H"  ;
    if (arc_index == 2442) return "H"  ;
    if (arc_index == 2464) return "E"  ;
    if (arc_index == 2469) return "E"  ;
    if (arc_index == 2470) return "E"  ;
    if (arc_index == 2472) return "E"  ;
    if (arc_index == 2473) return "H"  ;
    if (arc_index == 2474) return "W"  ;
    if (arc_index == 2475) return "W"  ;
    if (arc_index == 2477) return "W"  ;
    if (arc_index == 2480) return "W"  ;
    if (arc_index == 2483) return "W"  ;
    if (arc_index == 2485) return "W"  ;
    if (arc_index == 2567) return "E"  ;
    if (arc_index == 2576) return "E"  ;
    if (arc_index == 2589) return "H"  ;
    if (arc_index == 2597) return "H"  ;
    if (arc_index == 2674) return "H"  ;
    if (arc_index == 2678) return "H"  ;
    if (arc_index == 2692) return "H"  ;
    if (arc_index == 2702) return "H"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2739) return "W"  ;
    if (arc_index == 2760) return "W"  ;
    if (arc_index == 2761) return "W"  ;
    if (arc_index == 2765) return "W"  ;
    if (arc_index == 2770) return "W"  ;
    if (arc_index == 2792) return "W"  ;
    if (arc_index == 2800) return "W"  ;
    if (arc_index == 2801) return "W"  ;
    if (arc_index == 2809) return "W"  ;
    if (arc_index == 2823) return "H"  ;
    if (arc_index == 2834) return "W"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2842) return "E"  ;
    if (arc_index == 2854) return "E"  ;
    if (arc_index == 2856) return "E"  ;
    if (arc_index == 2861) return "E"  ;
    if (arc_index == 2893) return "E"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 5)) begin 
    if (arc_index == 28) return "E"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 72) return "H"  ;
    if (arc_index == 98) return "H"  ;
    if (arc_index == 130) return "H"  ;
    if (arc_index == 142) return "H"  ;
    if (arc_index == 216) return "H"  ;
    if (arc_index == 239) return "H"  ;
    if (arc_index == 333) return "H"  ;
    if (arc_index == 367) return "H"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 412) return "E"  ;
    if (arc_index == 414) return "E"  ;
    if (arc_index == 475) return "E"  ;
    if (arc_index == 480) return "E"  ;
    if (arc_index == 482) return "E"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 512) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 553) return "W"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 593) return "E"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 609) return "W"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 634) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 721) return "H"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 757) return "W"  ;
    if (arc_index == 759) return "W"  ;
    if (arc_index == 765) return "W"  ;
    if (arc_index == 784) return "W"  ;
    if (arc_index == 819) return "W"  ;
    if (arc_index == 822) return "W"  ;
    if (arc_index == 837) return "W"  ;
    if (arc_index == 876) return "H"  ;
    if (arc_index == 879) return "H"  ;
    if (arc_index == 882) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 965) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1009) return "H"  ;
    if (arc_index == 1017) return "H"  ;
    if (arc_index == 1056) return "W"  ;
    if (arc_index == 1078) return "E"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1092) return "E"  ;
    if (arc_index == 1093) return "E"  ;
    if (arc_index == 1104) return "H"  ;
    if (arc_index == 1105) return "W"  ;
    if (arc_index == 1106) return "W"  ;
    if (arc_index == 1110) return "W"  ;
    if (arc_index == 1111) return "W"  ;
    if (arc_index == 1121) return "W"  ;
    if (arc_index == 1149) return "W"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1190) return "E"  ;
    if (arc_index == 1230) return "H"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1341) return "H"  ;
    if (arc_index == 1344) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1390) return "W"  ;
    if (arc_index == 1393) return "W"  ;
    if (arc_index == 1397) return "W"  ;
    if (arc_index == 1408) return "W"  ;
    if (arc_index == 1411) return "H"  ;
    if (arc_index == 1428) return "W"  ;
    if (arc_index == 1430) return "W"  ;
    if (arc_index == 1432) return "W"  ;
    if (arc_index == 1441) return "W"  ;
    if (arc_index == 1453) return "W"  ;
    if (arc_index == 1455) return "W"  ;
    if (arc_index == 1463) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1498) return "W"  ;
    if (arc_index == 1514) return "W"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1541) return "W"  ;
    if (arc_index == 1586) return "H"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1610) return "E"  ;
    if (arc_index == 1613) return "E"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1619) return "E"  ;
    if (arc_index == 1620) return "E"  ;
    if (arc_index == 1624) return "E"  ;
    if (arc_index == 1638) return "E"  ;
    if (arc_index == 1650) return "E"  ;
    if (arc_index == 1653) return "E"  ;
    if (arc_index == 1654) return "E"  ;
    if (arc_index == 1666) return "E"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1672) return "E"  ;
    if (arc_index == 1673) return "W"  ;
    if (arc_index == 1691) return "W"  ;
    if (arc_index == 1696) return "W"  ;
    if (arc_index == 1698) return "W"  ;
    if (arc_index == 1707) return "W"  ;
    if (arc_index == 1710) return "W"  ;
    if (arc_index == 1730) return "W"  ;
    if (arc_index == 1734) return "W"  ;
    if (arc_index == 1737) return "E"  ;
    if (arc_index == 1747) return "E"  ;
    if (arc_index == 1773) return "E"  ;
    if (arc_index == 1776) return "E"  ;
    if (arc_index == 1783) return "H"  ;
    if (arc_index == 1789) return "H"  ;
    if (arc_index == 1790) return "W"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1802) return "W"  ;
    if (arc_index == 1804) return "W"  ;
    if (arc_index == 1812) return "W"  ;
    if (arc_index == 1822) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1826) return "H"  ;
    if (arc_index == 1829) return "E"  ;
    if (arc_index == 1848) return "E"  ;
    if (arc_index == 1849) return "W"  ;
    if (arc_index == 1850) return "W"  ;
    if (arc_index == 1851) return "E"  ;
    if (arc_index == 1852) return "E"  ;
    if (arc_index == 1853) return "W"  ;
    if (arc_index == 1854) return "W"  ;
    if (arc_index == 1855) return "W"  ;
    if (arc_index == 1856) return "W"  ;
    if (arc_index == 1857) return "W"  ;
    if (arc_index == 1858) return "E"  ;
    if (arc_index == 1859) return "E"  ;
    if (arc_index == 1860) return "E"  ;
    if (arc_index == 1861) return "W"  ;
    if (arc_index == 1862) return "W"  ;
    if (arc_index == 1863) return "E"  ;
    if (arc_index == 1864) return "E"  ;
    if (arc_index == 1865) return "E"  ;
    if (arc_index == 1866) return "E"  ;
    if (arc_index == 1867) return "E"  ;
    if (arc_index == 1868) return "E"  ;
    if (arc_index == 1869) return "E"  ;
    if (arc_index == 1877) return "E"  ;
    if (arc_index == 1881) return "H"  ;
    if (arc_index == 1889) return "H"  ;
    if (arc_index == 1892) return "W"  ;
    if (arc_index == 1895) return "W"  ;
    if (arc_index == 1898) return "W"  ;
    if (arc_index == 1904) return "W"  ;
    if (arc_index == 1906) return "E"  ;
    if (arc_index == 1911) return "W"  ;
    if (arc_index == 1912) return "W"  ;
    if (arc_index == 1917) return "E"  ;
    if (arc_index == 1924) return "E"  ;
    if (arc_index == 1925) return "E"  ;
    if (arc_index == 1926) return "H"  ;
    if (arc_index == 1928) return "E"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1952) return "E"  ;
    if (arc_index == 1982) return "E"  ;
    if (arc_index == 1988) return "E"  ;
    if (arc_index == 1994) return "E"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2049) return "E"  ;
    if (arc_index == 2059) return "E"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2091) return "W"  ;
    if (arc_index == 2115) return "W"  ;
    if (arc_index == 2121) return "E"  ;
    if (arc_index == 2123) return "E"  ;
    if (arc_index == 2125) return "H"  ;
    if (arc_index == 2132) return "W"  ;
    if (arc_index == 2152) return "E"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2188) return "W"  ;
    if (arc_index == 2202) return "W"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2224) return "W"  ;
    if (arc_index == 2238) return "W"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2254) return "W"  ;
    if (arc_index == 2257) return "W"  ;
    if (arc_index == 2280) return "W"  ;
    if (arc_index == 2302) return "H"  ;
    if (arc_index == 2313) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2363) return "W"  ;
    if (arc_index == 2368) return "W"  ;
    if (arc_index == 2369) return "W"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2375) return "W"  ;
    if (arc_index == 2386) return "H"  ;
    if (arc_index == 2413) return "W"  ;
    if (arc_index == 2421) return "W"  ;
    if (arc_index == 2424) return "E"  ;
    if (arc_index == 2429) return "E"  ;
    if (arc_index == 2486) return "W"  ;
    if (arc_index == 2489) return "W"  ;
    if (arc_index == 2491) return "W"  ;
    if (arc_index == 2493) return "W"  ;
    if (arc_index == 2494) return "W"  ;
    if (arc_index == 2495) return "H"  ;
    if (arc_index == 2498) return "H"  ;
    if (arc_index == 2499) return "W"  ;
    if (arc_index == 2500) return "W"  ;
    if (arc_index == 2505) return "W"  ;
    if (arc_index == 2507) return "E"  ;
    if (arc_index == 2519) return "E"  ;
    if (arc_index == 2533) return "E"  ;
    if (arc_index == 2534) return "E"  ;
    if (arc_index == 2535) return "E"  ;
    if (arc_index == 2537) return "E"  ;
    if (arc_index == 2539) return "E"  ;
    if (arc_index == 2540) return "W"  ;
    if (arc_index == 2541) return "W"  ;
    if (arc_index == 2549) return "W"  ;
    if (arc_index == 2551) return "W"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2603) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2611) return "H"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2627) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2687) return "E"  ;
    if (arc_index == 2700) return "H"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2707) return "E"  ;
    if (arc_index == 2714) return "H"  ;
    if (arc_index == 2736) return "H"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2744) return "E"  ;
    if (arc_index == 2749) return "E"  ;
    if (arc_index == 2758) return "E"  ;
    if (arc_index == 2759) return "E"  ;
    if (arc_index == 2764) return "E"  ;
    if (arc_index == 2767) return "E"  ;
    if (arc_index == 2771) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2801) return "E"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2817) return "W"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2841) return "E"  ;
    if (arc_index == 2845) return "H"  ;
    if (arc_index == 2847) return "H"  ;
    if (arc_index == 2882) return "H"  ;
    if (arc_index == 2892) return "E"  ;
    if (arc_index == 2899) return "E"  ;
    if (arc_index == 2919) return "E"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 8)) begin 
    if (arc_index == 24) return "W"  ;
    if (arc_index == 31) return "E"  ;
    if (arc_index == 62) return "E"  ;
    if (arc_index == 89) return "E"  ;
    if (arc_index == 94) return "H"  ;
    if (arc_index == 104) return "E"  ;
    if (arc_index == 111) return "E"  ;
    if (arc_index == 154) return "E"  ;
    if (arc_index == 163) return "W"  ;
    if (arc_index == 166) return "W"  ;
    if (arc_index == 171) return "W"  ;
    if (arc_index == 176) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 180) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 182) return "W"  ;
    if (arc_index == 184) return "W"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 187) return "W"  ;
    if (arc_index == 188) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 194) return "W"  ;
    if (arc_index == 219) return "W"  ;
    if (arc_index == 229) return "W"  ;
    if (arc_index == 237) return "W"  ;
    if (arc_index == 240) return "W"  ;
    if (arc_index == 252) return "W"  ;
    if (arc_index == 260) return "W"  ;
    if (arc_index == 271) return "W"  ;
    if (arc_index == 279) return "W"  ;
    if (arc_index == 282) return "W"  ;
    if (arc_index == 287) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 304) return "W"  ;
    if (arc_index == 364) return "W"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 420) return "E"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 531) return "W"  ;
    if (arc_index == 532) return "W"  ;
    if (arc_index == 542) return "W"  ;
    if (arc_index == 548) return "W"  ;
    if (arc_index == 554) return "W"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 596) return "E"  ;
    if (arc_index == 616) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 636) return "W"  ;
    if (arc_index == 646) return "E"  ;
    if (arc_index == 704) return "E"  ;
    if (arc_index == 730) return "E"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 736) return "W"  ;
    if (arc_index == 737) return "E"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 743) return "H"  ;
    if (arc_index == 791) return "H"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 817) return "E"  ;
    if (arc_index == 825) return "E"  ;
    if (arc_index == 867) return "E"  ;
    if (arc_index == 898) return "H"  ;
    if (arc_index == 933) return "H"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 969) return "E"  ;
    if (arc_index == 982) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1031) return "H"  ;
    if (arc_index == 1035) return "W"  ;
    if (arc_index == 1039) return "H"  ;
    if (arc_index == 1040) return "H"  ;
    if (arc_index == 1057) return "E"  ;
    if (arc_index == 1073) return "E"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1100) return "E"  ;
    if (arc_index == 1126) return "H"  ;
    if (arc_index == 1127) return "H"  ;
    if (arc_index == 1140) return "H"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1167) return "W"  ;
    if (arc_index == 1173) return "E"  ;
    if (arc_index == 1183) return "E"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1236) return "E"  ;
    if (arc_index == 1244) return "W"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1252) return "H"  ;
    if (arc_index == 1254) return "W"  ;
    if (arc_index == 1255) return "W"  ;
    if (arc_index == 1257) return "W"  ;
    if (arc_index == 1259) return "W"  ;
    if (arc_index == 1261) return "W"  ;
    if (arc_index == 1263) return "W"  ;
    if (arc_index == 1266) return "W"  ;
    if (arc_index == 1268) return "E"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1271) return "E"  ;
    if (arc_index == 1273) return "W"  ;
    if (arc_index == 1274) return "W"  ;
    if (arc_index == 1275) return "W"  ;
    if (arc_index == 1276) return "W"  ;
    if (arc_index == 1278) return "E"  ;
    if (arc_index == 1283) return "E"  ;
    if (arc_index == 1302) return "E"  ;
    if (arc_index == 1332) return "E"  ;
    if (arc_index == 1361) return "E"  ;
    if (arc_index == 1363) return "H"  ;
    if (arc_index == 1370) return "H"  ;
    if (arc_index == 1382) return "H"  ;
    if (arc_index == 1433) return "H"  ;
    if (arc_index == 1471) return "E"  ;
    if (arc_index == 1489) return "E"  ;
    if (arc_index == 1501) return "E"  ;
    if (arc_index == 1550) return "E"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1608) return "H"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1677) return "W"  ;
    if (arc_index == 1693) return "W"  ;
    if (arc_index == 1708) return "W"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1763) return "E"  ;
    if (arc_index == 1792) return "E"  ;
    if (arc_index == 1803) return "E"  ;
    if (arc_index == 1805) return "H"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1848) return "H"  ;
    if (arc_index == 1870) return "H"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1872) return "W"  ;
    if (arc_index == 1873) return "E"  ;
    if (arc_index == 1874) return "E"  ;
    if (arc_index == 1875) return "E"  ;
    if (arc_index == 1876) return "E"  ;
    if (arc_index == 1877) return "E"  ;
    if (arc_index == 1878) return "W"  ;
    if (arc_index == 1879) return "W"  ;
    if (arc_index == 1880) return "W"  ;
    if (arc_index == 1881) return "W"  ;
    if (arc_index == 1882) return "W"  ;
    if (arc_index == 1883) return "W"  ;
    if (arc_index == 1884) return "W"  ;
    if (arc_index == 1885) return "W"  ;
    if (arc_index == 1886) return "E"  ;
    if (arc_index == 1887) return "E"  ;
    if (arc_index == 1888) return "E"  ;
    if (arc_index == 1889) return "E"  ;
    if (arc_index == 1890) return "E"  ;
    if (arc_index == 1891) return "E"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 1900) return "E"  ;
    if (arc_index == 1901) return "E"  ;
    if (arc_index == 1903) return "H"  ;
    if (arc_index == 1938) return "H"  ;
    if (arc_index == 1948) return "H"  ;
    if (arc_index == 1995) return "H"  ;
    if (arc_index == 2019) return "H"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2077) return "W"  ;
    if (arc_index == 2087) return "W"  ;
    if (arc_index == 2106) return "W"  ;
    if (arc_index == 2130) return "E"  ;
    if (arc_index == 2133) return "E"  ;
    if (arc_index == 2136) return "E"  ;
    if (arc_index == 2147) return "H"  ;
    if (arc_index == 2183) return "H"  ;
    if (arc_index == 2206) return "W"  ;
    if (arc_index == 2210) return "W"  ;
    if (arc_index == 2214) return "W"  ;
    if (arc_index == 2215) return "W"  ;
    if (arc_index == 2218) return "W"  ;
    if (arc_index == 2263) return "E"  ;
    if (arc_index == 2272) return "E"  ;
    if (arc_index == 2278) return "E"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2314) return "W"  ;
    if (arc_index == 2316) return "W"  ;
    if (arc_index == 2318) return "W"  ;
    if (arc_index == 2319) return "W"  ;
    if (arc_index == 2321) return "W"  ;
    if (arc_index == 2323) return "W"  ;
    if (arc_index == 2324) return "H"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2330) return "W"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2361) return "W"  ;
    if (arc_index == 2404) return "W"  ;
    if (arc_index == 2408) return "H"  ;
    if (arc_index == 2411) return "H"  ;
    if (arc_index == 2444) return "E"  ;
    if (arc_index == 2462) return "E"  ;
    if (arc_index == 2517) return "H"  ;
    if (arc_index == 2528) return "H"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2599) return "W"  ;
    if (arc_index == 2600) return "W"  ;
    if (arc_index == 2633) return "H"  ;
    if (arc_index == 2644) return "H"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2719) return "E"  ;
    if (arc_index == 2722) return "H"  ;
    if (arc_index == 2725) return "W"  ;
    if (arc_index == 2736) return "H"  ;
    if (arc_index == 2738) return "H"  ;
    if (arc_index == 2764) return "E"  ;
    if (arc_index == 2821) return "E"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2867) return "H"  ;
    if (arc_index == 2907) return "H"  ;
    if (arc_index == 2908) return "H"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 5)) begin 
    if (arc_index == 0) return "H"  ;
    if (arc_index == 7) return "W"  ;
    if (arc_index == 13) return "W"  ;
    if (arc_index == 18) return "W"  ;
    if (arc_index == 30) return "E"  ;
    if (arc_index == 72) return "E"  ;
    if (arc_index == 78) return "E"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 98) return "E"  ;
    if (arc_index == 101) return "W"  ;
    if (arc_index == 116) return "H"  ;
    if (arc_index == 130) return "H"  ;
    if (arc_index == 142) return "H"  ;
    if (arc_index == 158) return "W"  ;
    if (arc_index == 159) return "W"  ;
    if (arc_index == 160) return "W"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 212) return "W"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 233) return "W"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 296) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 367) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 386) return "W"  ;
    if (arc_index == 399) return "E"  ;
    if (arc_index == 412) return "E"  ;
    if (arc_index == 414) return "E"  ;
    if (arc_index == 454) return "E"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 535) return "W"  ;
    if (arc_index == 553) return "W"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 603) return "W"  ;
    if (arc_index == 609) return "W"  ;
    if (arc_index == 610) return "W"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 654) return "W"  ;
    if (arc_index == 663) return "E"  ;
    if (arc_index == 686) return "E"  ;
    if (arc_index == 687) return "E"  ;
    if (arc_index == 744) return "E"  ;
    if (arc_index == 757) return "E"  ;
    if (arc_index == 759) return "E"  ;
    if (arc_index == 765) return "H"  ;
    if (arc_index == 769) return "H"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 784) return "E"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 837) return "E"  ;
    if (arc_index == 876) return "E"  ;
    if (arc_index == 879) return "E"  ;
    if (arc_index == 898) return "E"  ;
    if (arc_index == 917) return "E"  ;
    if (arc_index == 920) return "H"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 971) return "E"  ;
    if (arc_index == 974) return "W"  ;
    if (arc_index == 1009) return "W"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1017) return "E"  ;
    if (arc_index == 1053) return "H"  ;
    if (arc_index == 1061) return "H"  ;
    if (arc_index == 1063) return "W"  ;
    if (arc_index == 1068) return "W"  ;
    if (arc_index == 1075) return "W"  ;
    if (arc_index == 1077) return "W"  ;
    if (arc_index == 1085) return "E"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1092) return "E"  ;
    if (arc_index == 1093) return "E"  ;
    if (arc_index == 1106) return "W"  ;
    if (arc_index == 1121) return "W"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1148) return "H"  ;
    if (arc_index == 1170) return "W"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1230) return "E"  ;
    if (arc_index == 1274) return "H"  ;
    if (arc_index == 1279) return "W"  ;
    if (arc_index == 1280) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1385) return "H"  ;
    if (arc_index == 1393) return "H"  ;
    if (arc_index == 1397) return "E"  ;
    if (arc_index == 1408) return "E"  ;
    if (arc_index == 1422) return "E"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1430) return "W"  ;
    if (arc_index == 1432) return "W"  ;
    if (arc_index == 1441) return "W"  ;
    if (arc_index == 1455) return "H"  ;
    if (arc_index == 1463) return "H"  ;
    if (arc_index == 1494) return "H"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1498) return "W"  ;
    if (arc_index == 1514) return "W"  ;
    if (arc_index == 1520) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1594) return "E"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1607) return "E"  ;
    if (arc_index == 1608) return "E"  ;
    if (arc_index == 1615) return "E"  ;
    if (arc_index == 1621) return "E"  ;
    if (arc_index == 1626) return "E"  ;
    if (arc_index == 1630) return "H"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1635) return "E"  ;
    if (arc_index == 1641) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1672) return "E"  ;
    if (arc_index == 1673) return "E"  ;
    if (arc_index == 1684) return "W"  ;
    if (arc_index == 1696) return "E"  ;
    if (arc_index == 1698) return "E"  ;
    if (arc_index == 1707) return "E"  ;
    if (arc_index == 1710) return "E"  ;
    if (arc_index == 1730) return "E"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1773) return "E"  ;
    if (arc_index == 1775) return "E"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1785) return "W"  ;
    if (arc_index == 1789) return "W"  ;
    if (arc_index == 1802) return "W"  ;
    if (arc_index == 1823) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1827) return "H"  ;
    if (arc_index == 1850) return "H"  ;
    if (arc_index == 1855) return "H"  ;
    if (arc_index == 1856) return "H"  ;
    if (arc_index == 1864) return "H"  ;
    if (arc_index == 1865) return "H"  ;
    if (arc_index == 1870) return "H"  ;
    if (arc_index == 1881) return "H"  ;
    if (arc_index == 1892) return "H"  ;
    if (arc_index == 1893) return "E"  ;
    if (arc_index == 1894) return "W"  ;
    if (arc_index == 1895) return "W"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 1897) return "W"  ;
    if (arc_index == 1898) return "W"  ;
    if (arc_index == 1899) return "W"  ;
    if (arc_index == 1900) return "W"  ;
    if (arc_index == 1901) return "E"  ;
    if (arc_index == 1902) return "E"  ;
    if (arc_index == 1903) return "E"  ;
    if (arc_index == 1904) return "E"  ;
    if (arc_index == 1905) return "W"  ;
    if (arc_index == 1906) return "W"  ;
    if (arc_index == 1907) return "E"  ;
    if (arc_index == 1908) return "E"  ;
    if (arc_index == 1909) return "E"  ;
    if (arc_index == 1910) return "W"  ;
    if (arc_index == 1911) return "W"  ;
    if (arc_index == 1912) return "W"  ;
    if (arc_index == 1913) return "W"  ;
    if (arc_index == 1916) return "W"  ;
    if (arc_index == 1922) return "E"  ;
    if (arc_index == 1925) return "H"  ;
    if (arc_index == 1936) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1953) return "E"  ;
    if (arc_index == 1954) return "E"  ;
    if (arc_index == 1969) return "W"  ;
    if (arc_index == 1970) return "H"  ;
    if (arc_index == 1982) return "E"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2032) return "E"  ;
    if (arc_index == 2036) return "E"  ;
    if (arc_index == 2042) return "E"  ;
    if (arc_index == 2049) return "E"  ;
    if (arc_index == 2053) return "E"  ;
    if (arc_index == 2059) return "E"  ;
    if (arc_index == 2090) return "E"  ;
    if (arc_index == 2091) return "E"  ;
    if (arc_index == 2115) return "E"  ;
    if (arc_index == 2121) return "E"  ;
    if (arc_index == 2122) return "W"  ;
    if (arc_index == 2123) return "W"  ;
    if (arc_index == 2125) return "W"  ;
    if (arc_index == 2132) return "W"  ;
    if (arc_index == 2160) return "W"  ;
    if (arc_index == 2169) return "H"  ;
    if (arc_index == 2188) return "H"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2202) return "W"  ;
    if (arc_index == 2237) return "E"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2247) return "W"  ;
    if (arc_index == 2253) return "W"  ;
    if (arc_index == 2254) return "W"  ;
    if (arc_index == 2264) return "W"  ;
    if (arc_index == 2276) return "W"  ;
    if (arc_index == 2346) return "H"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2421) return "W"  ;
    if (arc_index == 2424) return "W"  ;
    if (arc_index == 2429) return "W"  ;
    if (arc_index == 2430) return "H"  ;
    if (arc_index == 2449) return "E"  ;
    if (arc_index == 2489) return "E"  ;
    if (arc_index == 2491) return "E"  ;
    if (arc_index == 2493) return "E"  ;
    if (arc_index == 2498) return "E"  ;
    if (arc_index == 2500) return "E"  ;
    if (arc_index == 2505) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2533) return "E"  ;
    if (arc_index == 2534) return "E"  ;
    if (arc_index == 2535) return "W"  ;
    if (arc_index == 2537) return "E"  ;
    if (arc_index == 2539) return "H"  ;
    if (arc_index == 2541) return "W"  ;
    if (arc_index == 2549) return "W"  ;
    if (arc_index == 2551) return "W"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2620) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2655) return "H"  ;
    if (arc_index == 2664) return "E"  ;
    if (arc_index == 2670) return "E"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2687) return "E"  ;
    if (arc_index == 2689) return "E"  ;
    if (arc_index == 2690) return "E"  ;
    if (arc_index == 2696) return "E"  ;
    if (arc_index == 2698) return "E"  ;
    if (arc_index == 2700) return "E"  ;
    if (arc_index == 2705) return "E"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2736) return "W"  ;
    if (arc_index == 2739) return "W"  ;
    if (arc_index == 2744) return "H"  ;
    if (arc_index == 2758) return "H"  ;
    if (arc_index == 2759) return "H"  ;
    if (arc_index == 2764) return "H"  ;
    if (arc_index == 2767) return "H"  ;
    if (arc_index == 2771) return "H"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2841) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2861) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2889) return "H"  ;
    if (arc_index == 2894) return "E"  ;
    if (arc_index == 2895) return "E"  ;
    if (arc_index == 2902) return "E"  ;
    if (arc_index == 2912) return "E"  ;
    if (arc_index == 2915) return "W"  ;
    if (arc_index == 2919) return "W"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 2)) begin 
    if (arc_index == 65) return "W"  ;
    if (arc_index == 80) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 115) return "W"  ;
    if (arc_index == 136) return "W"  ;
    if (arc_index == 138) return "H"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 384) return "E"  ;
    if (arc_index == 390) return "E"  ;
    if (arc_index == 439) return "E"  ;
    if (arc_index == 443) return "E"  ;
    if (arc_index == 478) return "W"  ;
    if (arc_index == 485) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 512) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 521) return "E"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 523) return "E"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 574) return "E"  ;
    if (arc_index == 576) return "E"  ;
    if (arc_index == 578) return "E"  ;
    if (arc_index == 589) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 593) return "E"  ;
    if (arc_index == 605) return "W"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 654) return "W"  ;
    if (arc_index == 668) return "W"  ;
    if (arc_index == 751) return "W"  ;
    if (arc_index == 770) return "W"  ;
    if (arc_index == 779) return "W"  ;
    if (arc_index == 787) return "H"  ;
    if (arc_index == 789) return "H"  ;
    if (arc_index == 799) return "H"  ;
    if (arc_index == 803) return "H"  ;
    if (arc_index == 840) return "W"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 880) return "W"  ;
    if (arc_index == 884) return "W"  ;
    if (arc_index == 886) return "W"  ;
    if (arc_index == 888) return "W"  ;
    if (arc_index == 896) return "W"  ;
    if (arc_index == 898) return "E"  ;
    if (arc_index == 900) return "E"  ;
    if (arc_index == 906) return "E"  ;
    if (arc_index == 907) return "E"  ;
    if (arc_index == 909) return "E"  ;
    if (arc_index == 913) return "E"  ;
    if (arc_index == 931) return "E"  ;
    if (arc_index == 942) return "H"  ;
    if (arc_index == 953) return "H"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 965) return "E"  ;
    if (arc_index == 994) return "E"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1056) return "W"  ;
    if (arc_index == 1075) return "H"  ;
    if (arc_index == 1083) return "H"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1099) return "E"  ;
    if (arc_index == 1105) return "E"  ;
    if (arc_index == 1110) return "W"  ;
    if (arc_index == 1111) return "W"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1170) return "H"  ;
    if (arc_index == 1193) return "H"  ;
    if (arc_index == 1202) return "H"  ;
    if (arc_index == 1209) return "H"  ;
    if (arc_index == 1213) return "E"  ;
    if (arc_index == 1231) return "E"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1296) return "H"  ;
    if (arc_index == 1335) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1391) return "W"  ;
    if (arc_index == 1407) return "H"  ;
    if (arc_index == 1438) return "W"  ;
    if (arc_index == 1453) return "W"  ;
    if (arc_index == 1477) return "H"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1527) return "W"  ;
    if (arc_index == 1533) return "W"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1584) return "E"  ;
    if (arc_index == 1585) return "E"  ;
    if (arc_index == 1586) return "E"  ;
    if (arc_index == 1587) return "E"  ;
    if (arc_index == 1588) return "E"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1616) return "E"  ;
    if (arc_index == 1628) return "E"  ;
    if (arc_index == 1636) return "E"  ;
    if (arc_index == 1643) return "E"  ;
    if (arc_index == 1647) return "E"  ;
    if (arc_index == 1652) return "H"  ;
    if (arc_index == 1656) return "W"  ;
    if (arc_index == 1661) return "W"  ;
    if (arc_index == 1662) return "W"  ;
    if (arc_index == 1664) return "W"  ;
    if (arc_index == 1665) return "W"  ;
    if (arc_index == 1673) return "W"  ;
    if (arc_index == 1706) return "W"  ;
    if (arc_index == 1719) return "W"  ;
    if (arc_index == 1723) return "W"  ;
    if (arc_index == 1726) return "W"  ;
    if (arc_index == 1731) return "W"  ;
    if (arc_index == 1735) return "W"  ;
    if (arc_index == 1740) return "W"  ;
    if (arc_index == 1743) return "W"  ;
    if (arc_index == 1752) return "W"  ;
    if (arc_index == 1754) return "W"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1830) return "W"  ;
    if (arc_index == 1831) return "W"  ;
    if (arc_index == 1849) return "H"  ;
    if (arc_index == 1861) return "W"  ;
    if (arc_index == 1892) return "H"  ;
    if (arc_index == 1897) return "H"  ;
    if (arc_index == 1914) return "H"  ;
    if (arc_index == 1915) return "H"  ;
    if (arc_index == 1916) return "E"  ;
    if (arc_index == 1917) return "E"  ;
    if (arc_index == 1918) return "W"  ;
    if (arc_index == 1919) return "W"  ;
    if (arc_index == 1920) return "W"  ;
    if (arc_index == 1921) return "W"  ;
    if (arc_index == 1922) return "E"  ;
    if (arc_index == 1923) return "E"  ;
    if (arc_index == 1924) return "E"  ;
    if (arc_index == 1925) return "E"  ;
    if (arc_index == 1926) return "E"  ;
    if (arc_index == 1927) return "E"  ;
    if (arc_index == 1928) return "E"  ;
    if (arc_index == 1929) return "E"  ;
    if (arc_index == 1930) return "W"  ;
    if (arc_index == 1931) return "W"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1933) return "E"  ;
    if (arc_index == 1934) return "E"  ;
    if (arc_index == 1935) return "E"  ;
    if (arc_index == 1941) return "E"  ;
    if (arc_index == 1947) return "H"  ;
    if (arc_index == 1992) return "H"  ;
    if (arc_index == 2002) return "H"  ;
    if (arc_index == 2007) return "E"  ;
    if (arc_index == 2015) return "E"  ;
    if (arc_index == 2115) return "W"  ;
    if (arc_index == 2191) return "H"  ;
    if (arc_index == 2223) return "E"  ;
    if (arc_index == 2238) return "E"  ;
    if (arc_index == 2368) return "H"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2452) return "H"  ;
    if (arc_index == 2460) return "W"  ;
    if (arc_index == 2480) return "W"  ;
    if (arc_index == 2494) return "W"  ;
    if (arc_index == 2499) return "W"  ;
    if (arc_index == 2526) return "W"  ;
    if (arc_index == 2555) return "W"  ;
    if (arc_index == 2557) return "E"  ;
    if (arc_index == 2561) return "H"  ;
    if (arc_index == 2566) return "H"  ;
    if (arc_index == 2576) return "H"  ;
    if (arc_index == 2582) return "H"  ;
    if (arc_index == 2590) return "H"  ;
    if (arc_index == 2597) return "H"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2674) return "W"  ;
    if (arc_index == 2677) return "H"  ;
    if (arc_index == 2678) return "E"  ;
    if (arc_index == 2679) return "E"  ;
    if (arc_index == 2688) return "W"  ;
    if (arc_index == 2733) return "W"  ;
    if (arc_index == 2754) return "W"  ;
    if (arc_index == 2760) return "W"  ;
    if (arc_index == 2765) return "W"  ;
    if (arc_index == 2766) return "H"  ;
    if (arc_index == 2778) return "H"  ;
    if (arc_index == 2780) return "H"  ;
    if (arc_index == 2788) return "H"  ;
    if (arc_index == 2803) return "E"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2812) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2868) return "E"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2881) return "E"  ;
    if (arc_index == 2900) return "E"  ;
    if (arc_index == 2911) return "H"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 1)) begin 
    if (arc_index == 7) return "H"  ;
    if (arc_index == 69) return "H"  ;
    if (arc_index == 79) return "H"  ;
    if (arc_index == 106) return "H"  ;
    if (arc_index == 145) return "H"  ;
    if (arc_index == 160) return "H"  ;
    if (arc_index == 384) return "E"  ;
    if (arc_index == 389) return "E"  ;
    if (arc_index == 406) return "E"  ;
    if (arc_index == 441) return "E"  ;
    if (arc_index == 449) return "E"  ;
    if (arc_index == 450) return "E"  ;
    if (arc_index == 460) return "E"  ;
    if (arc_index == 484) return "E"  ;
    if (arc_index == 486) return "E"  ;
    if (arc_index == 494) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 513) return "E"  ;
    if (arc_index == 514) return "E"  ;
    if (arc_index == 517) return "E"  ;
    if (arc_index == 518) return "E"  ;
    if (arc_index == 520) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 591) return "E"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 641) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 773) return "W"  ;
    if (arc_index == 774) return "W"  ;
    if (arc_index == 800) return "W"  ;
    if (arc_index == 809) return "H"  ;
    if (arc_index == 894) return "H"  ;
    if (arc_index == 924) return "H"  ;
    if (arc_index == 946) return "E"  ;
    if (arc_index == 948) return "E"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 964) return "H"  ;
    if (arc_index == 979) return "H"  ;
    if (arc_index == 1013) return "H"  ;
    if (arc_index == 1018) return "H"  ;
    if (arc_index == 1024) return "H"  ;
    if (arc_index == 1077) return "W"  ;
    if (arc_index == 1081) return "W"  ;
    if (arc_index == 1087) return "W"  ;
    if (arc_index == 1090) return "W"  ;
    if (arc_index == 1095) return "W"  ;
    if (arc_index == 1097) return "H"  ;
    if (arc_index == 1105) return "H"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1192) return "H"  ;
    if (arc_index == 1223) return "H"  ;
    if (arc_index == 1224) return "H"  ;
    if (arc_index == 1318) return "H"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1391) return "W"  ;
    if (arc_index == 1429) return "H"  ;
    if (arc_index == 1453) return "W"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1499) return "H"  ;
    if (arc_index == 1532) return "H"  ;
    if (arc_index == 1534) return "H"  ;
    if (arc_index == 1584) return "E"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1594) return "E"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1599) return "E"  ;
    if (arc_index == 1604) return "E"  ;
    if (arc_index == 1605) return "E"  ;
    if (arc_index == 1617) return "W"  ;
    if (arc_index == 1674) return "H"  ;
    if (arc_index == 1748) return "H"  ;
    if (arc_index == 1830) return "H"  ;
    if (arc_index == 1871) return "H"  ;
    if (arc_index == 1914) return "H"  ;
    if (arc_index == 1918) return "W"  ;
    if (arc_index == 1936) return "E"  ;
    if (arc_index == 1937) return "E"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1940) return "E"  ;
    if (arc_index == 1941) return "E"  ;
    if (arc_index == 1942) return "E"  ;
    if (arc_index == 1943) return "E"  ;
    if (arc_index == 1944) return "E"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1946) return "E"  ;
    if (arc_index == 1947) return "E"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1949) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 1951) return "E"  ;
    if (arc_index == 1952) return "E"  ;
    if (arc_index == 1953) return "E"  ;
    if (arc_index == 1954) return "E"  ;
    if (arc_index == 1955) return "E"  ;
    if (arc_index == 1956) return "E"  ;
    if (arc_index == 1957) return "E"  ;
    if (arc_index == 1969) return "H"  ;
    if (arc_index == 2014) return "H"  ;
    if (arc_index == 2021) return "W"  ;
    if (arc_index == 2116) return "W"  ;
    if (arc_index == 2122) return "W"  ;
    if (arc_index == 2176) return "W"  ;
    if (arc_index == 2213) return "H"  ;
    if (arc_index == 2221) return "H"  ;
    if (arc_index == 2223) return "E"  ;
    if (arc_index == 2224) return "E"  ;
    if (arc_index == 2228) return "E"  ;
    if (arc_index == 2232) return "E"  ;
    if (arc_index == 2238) return "E"  ;
    if (arc_index == 2242) return "E"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2390) return "H"  ;
    if (arc_index == 2423) return "W"  ;
    if (arc_index == 2450) return "W"  ;
    if (arc_index == 2474) return "H"  ;
    if (arc_index == 2499) return "H"  ;
    if (arc_index == 2552) return "H"  ;
    if (arc_index == 2556) return "H"  ;
    if (arc_index == 2571) return "W"  ;
    if (arc_index == 2582) return "E"  ;
    if (arc_index == 2583) return "H"  ;
    if (arc_index == 2585) return "H"  ;
    if (arc_index == 2593) return "H"  ;
    if (arc_index == 2607) return "H"  ;
    if (arc_index == 2670) return "E"  ;
    if (arc_index == 2695) return "W"  ;
    if (arc_index == 2699) return "H"  ;
    if (arc_index == 2730) return "H"  ;
    if (arc_index == 2746) return "E"  ;
    if (arc_index == 2747) return "E"  ;
    if (arc_index == 2748) return "E"  ;
    if (arc_index == 2760) return "E"  ;
    if (arc_index == 2788) return "H"  ;
    if (arc_index == 2796) return "H"  ;
    if (arc_index == 2802) return "H"  ;
    if (arc_index == 2811) return "H"  ;
    if (arc_index == 2851) return "H"  ;
    if (arc_index == 2859) return "H"  ;
    if (arc_index == 2860) return "E"  ;
    if (arc_index == 2863) return "E"  ;
    if (arc_index == 2869) return "E"  ;
    if (arc_index == 2903) return "W"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 7)) begin 
    if (arc_index == 21) return "W"  ;
    if (arc_index == 29) return "H"  ;
    if (arc_index == 43) return "H"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 92) return "E"  ;
    if (arc_index == 95) return "E"  ;
    if (arc_index == 97) return "E"  ;
    if (arc_index == 101) return "W"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 156) return "E"  ;
    if (arc_index == 165) return "E"  ;
    if (arc_index == 174) return "E"  ;
    if (arc_index == 176) return "E"  ;
    if (arc_index == 182) return "H"  ;
    if (arc_index == 183) return "W"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 201) return "W"  ;
    if (arc_index == 206) return "W"  ;
    if (arc_index == 233) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 270) return "W"  ;
    if (arc_index == 284) return "W"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 338) return "E"  ;
    if (arc_index == 342) return "E"  ;
    if (arc_index == 347) return "E"  ;
    if (arc_index == 354) return "E"  ;
    if (arc_index == 359) return "E"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 428) return "E"  ;
    if (arc_index == 431) return "E"  ;
    if (arc_index == 433) return "E"  ;
    if (arc_index == 438) return "E"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 463) return "E"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 469) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 481) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 535) return "W"  ;
    if (arc_index == 537) return "W"  ;
    if (arc_index == 539) return "W"  ;
    if (arc_index == 554) return "E"  ;
    if (arc_index == 561) return "E"  ;
    if (arc_index == 564) return "W"  ;
    if (arc_index == 595) return "W"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 607) return "W"  ;
    if (arc_index == 643) return "W"  ;
    if (arc_index == 652) return "W"  ;
    if (arc_index == 677) return "W"  ;
    if (arc_index == 695) return "W"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 736) return "W"  ;
    if (arc_index == 742) return "W"  ;
    if (arc_index == 772) return "W"  ;
    if (arc_index == 777) return "W"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 828) return "E"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 831) return "H"  ;
    if (arc_index == 857) return "H"  ;
    if (arc_index == 911) return "E"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 928) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 973) return "E"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 986) return "H"  ;
    if (arc_index == 1020) return "H"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1035) return "E"  ;
    if (arc_index == 1053) return "W"  ;
    if (arc_index == 1057) return "W"  ;
    if (arc_index == 1059) return "W"  ;
    if (arc_index == 1065) return "W"  ;
    if (arc_index == 1069) return "W"  ;
    if (arc_index == 1072) return "W"  ;
    if (arc_index == 1073) return "E"  ;
    if (arc_index == 1074) return "W"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1112) return "E"  ;
    if (arc_index == 1119) return "H"  ;
    if (arc_index == 1124) return "W"  ;
    if (arc_index == 1127) return "H"  ;
    if (arc_index == 1140) return "W"  ;
    if (arc_index == 1144) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1177) return "W"  ;
    if (arc_index == 1186) return "W"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1214) return "H"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1273) return "W"  ;
    if (arc_index == 1274) return "W"  ;
    if (arc_index == 1275) return "W"  ;
    if (arc_index == 1277) return "E"  ;
    if (arc_index == 1280) return "E"  ;
    if (arc_index == 1286) return "E"  ;
    if (arc_index == 1290) return "E"  ;
    if (arc_index == 1297) return "E"  ;
    if (arc_index == 1302) return "W"  ;
    if (arc_index == 1313) return "W"  ;
    if (arc_index == 1325) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1340) return "H"  ;
    if (arc_index == 1354) return "H"  ;
    if (arc_index == 1364) return "H"  ;
    if (arc_index == 1367) return "H"  ;
    if (arc_index == 1374) return "H"  ;
    if (arc_index == 1375) return "H"  ;
    if (arc_index == 1379) return "H"  ;
    if (arc_index == 1427) return "H"  ;
    if (arc_index == 1445) return "H"  ;
    if (arc_index == 1451) return "H"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1490) return "W"  ;
    if (arc_index == 1510) return "W"  ;
    if (arc_index == 1515) return "W"  ;
    if (arc_index == 1521) return "H"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1541) return "E"  ;
    if (arc_index == 1542) return "E"  ;
    if (arc_index == 1543) return "E"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1607) return "E"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1650) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1674) return "W"  ;
    if (arc_index == 1675) return "W"  ;
    if (arc_index == 1676) return "W"  ;
    if (arc_index == 1683) return "W"  ;
    if (arc_index == 1684) return "W"  ;
    if (arc_index == 1687) return "W"  ;
    if (arc_index == 1690) return "W"  ;
    if (arc_index == 1691) return "W"  ;
    if (arc_index == 1696) return "H"  ;
    if (arc_index == 1730) return "H"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1764) return "E"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1803) return "E"  ;
    if (arc_index == 1810) return "E"  ;
    if (arc_index == 1813) return "W"  ;
    if (arc_index == 1814) return "W"  ;
    if (arc_index == 1818) return "W"  ;
    if (arc_index == 1820) return "W"  ;
    if (arc_index == 1821) return "W"  ;
    if (arc_index == 1829) return "W"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1870) return "W"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1893) return "H"  ;
    if (arc_index == 1901) return "E"  ;
    if (arc_index == 1936) return "H"  ;
    if (arc_index == 1949) return "E"  ;
    if (arc_index == 1958) return "E"  ;
    if (arc_index == 1959) return "E"  ;
    if (arc_index == 1960) return "W"  ;
    if (arc_index == 1961) return "E"  ;
    if (arc_index == 1962) return "E"  ;
    if (arc_index == 1963) return "E"  ;
    if (arc_index == 1964) return "E"  ;
    if (arc_index == 1965) return "W"  ;
    if (arc_index == 1966) return "W"  ;
    if (arc_index == 1967) return "E"  ;
    if (arc_index == 1968) return "W"  ;
    if (arc_index == 1969) return "W"  ;
    if (arc_index == 1970) return "W"  ;
    if (arc_index == 1971) return "W"  ;
    if (arc_index == 1972) return "W"  ;
    if (arc_index == 1973) return "W"  ;
    if (arc_index == 1974) return "E"  ;
    if (arc_index == 1975) return "E"  ;
    if (arc_index == 1976) return "E"  ;
    if (arc_index == 1977) return "E"  ;
    if (arc_index == 1978) return "E"  ;
    if (arc_index == 1979) return "E"  ;
    if (arc_index == 1991) return "H"  ;
    if (arc_index == 1994) return "E"  ;
    if (arc_index == 2036) return "H"  ;
    if (arc_index == 2042) return "H"  ;
    if (arc_index == 2046) return "H"  ;
    if (arc_index == 2063) return "E"  ;
    if (arc_index == 2079) return "W"  ;
    if (arc_index == 2087) return "W"  ;
    if (arc_index == 2114) return "E"  ;
    if (arc_index == 2126) return "E"  ;
    if (arc_index == 2172) return "E"  ;
    if (arc_index == 2188) return "W"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2206) return "W"  ;
    if (arc_index == 2235) return "H"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2244) return "E"  ;
    if (arc_index == 2266) return "E"  ;
    if (arc_index == 2268) return "E"  ;
    if (arc_index == 2285) return "E"  ;
    if (arc_index == 2286) return "E"  ;
    if (arc_index == 2287) return "E"  ;
    if (arc_index == 2288) return "E"  ;
    if (arc_index == 2296) return "E"  ;
    if (arc_index == 2299) return "E"  ;
    if (arc_index == 2306) return "E"  ;
    if (arc_index == 2318) return "E"  ;
    if (arc_index == 2321) return "E"  ;
    if (arc_index == 2322) return "W"  ;
    if (arc_index == 2323) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2372) return "W"  ;
    if (arc_index == 2389) return "W"  ;
    if (arc_index == 2398) return "W"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2412) return "H"  ;
    if (arc_index == 2416) return "W"  ;
    if (arc_index == 2432) return "W"  ;
    if (arc_index == 2446) return "E"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2496) return "H"  ;
    if (arc_index == 2507) return "H"  ;
    if (arc_index == 2543) return "H"  ;
    if (arc_index == 2559) return "H"  ;
    if (arc_index == 2605) return "H"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2669) return "E"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2705) return "E"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2714) return "W"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2721) return "H"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2810) return "H"  ;
    if (arc_index == 2819) return "W"  ;
    if (arc_index == 2820) return "W"  ;
    if (arc_index == 2821) return "W"  ;
    if (arc_index == 2824) return "H"  ;
    if (arc_index == 2837) return "H"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2922) return "E"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 4)) begin 
    if (arc_index == 12) return "W"  ;
    if (arc_index == 51) return "H"  ;
    if (arc_index == 58) return "E"  ;
    if (arc_index == 86) return "E"  ;
    if (arc_index == 123) return "E"  ;
    if (arc_index == 130) return "E"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 200) return "W"  ;
    if (arc_index == 204) return "H"  ;
    if (arc_index == 211) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 244) return "W"  ;
    if (arc_index == 262) return "W"  ;
    if (arc_index == 301) return "W"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 384) return "W"  ;
    if (arc_index == 456) return "E"  ;
    if (arc_index == 470) return "E"  ;
    if (arc_index == 535) return "W"  ;
    if (arc_index == 550) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 571) return "W"  ;
    if (arc_index == 574) return "E"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 609) return "E"  ;
    if (arc_index == 611) return "E"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 688) return "W"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 699) return "W"  ;
    if (arc_index == 726) return "W"  ;
    if (arc_index == 750) return "W"  ;
    if (arc_index == 752) return "W"  ;
    if (arc_index == 754) return "E"  ;
    if (arc_index == 755) return "E"  ;
    if (arc_index == 756) return "E"  ;
    if (arc_index == 757) return "E"  ;
    if (arc_index == 758) return "E"  ;
    if (arc_index == 759) return "E"  ;
    if (arc_index == 761) return "E"  ;
    if (arc_index == 767) return "E"  ;
    if (arc_index == 769) return "E"  ;
    if (arc_index == 771) return "E"  ;
    if (arc_index == 775) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 784) return "E"  ;
    if (arc_index == 815) return "W"  ;
    if (arc_index == 840) return "W"  ;
    if (arc_index == 848) return "W"  ;
    if (arc_index == 849) return "W"  ;
    if (arc_index == 853) return "H"  ;
    if (arc_index == 854) return "W"  ;
    if (arc_index == 883) return "W"  ;
    if (arc_index == 887) return "E"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 892) return "E"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 901) return "E"  ;
    if (arc_index == 914) return "E"  ;
    if (arc_index == 949) return "E"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 961) return "E"  ;
    if (arc_index == 996) return "E"  ;
    if (arc_index == 1008) return "H"  ;
    if (arc_index == 1025) return "H"  ;
    if (arc_index == 1047) return "H"  ;
    if (arc_index == 1052) return "H"  ;
    if (arc_index == 1062) return "H"  ;
    if (arc_index == 1094) return "E"  ;
    if (arc_index == 1141) return "H"  ;
    if (arc_index == 1149) return "H"  ;
    if (arc_index == 1185) return "W"  ;
    if (arc_index == 1197) return "W"  ;
    if (arc_index == 1236) return "H"  ;
    if (arc_index == 1280) return "W"  ;
    if (arc_index == 1334) return "W"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1362) return "H"  ;
    if (arc_index == 1388) return "H"  ;
    if (arc_index == 1391) return "H"  ;
    if (arc_index == 1407) return "W"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1459) return "W"  ;
    if (arc_index == 1465) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1473) return "H"  ;
    if (arc_index == 1476) return "H"  ;
    if (arc_index == 1492) return "W"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1543) return "H"  ;
    if (arc_index == 1599) return "E"  ;
    if (arc_index == 1614) return "E"  ;
    if (arc_index == 1625) return "W"  ;
    if (arc_index == 1645) return "W"  ;
    if (arc_index == 1663) return "W"  ;
    if (arc_index == 1694) return "W"  ;
    if (arc_index == 1697) return "W"  ;
    if (arc_index == 1715) return "W"  ;
    if (arc_index == 1718) return "H"  ;
    if (arc_index == 1727) return "H"  ;
    if (arc_index == 1729) return "E"  ;
    if (arc_index == 1739) return "E"  ;
    if (arc_index == 1742) return "E"  ;
    if (arc_index == 1747) return "E"  ;
    if (arc_index == 1751) return "E"  ;
    if (arc_index == 1755) return "E"  ;
    if (arc_index == 1761) return "W"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1828) return "E"  ;
    if (arc_index == 1888) return "E"  ;
    if (arc_index == 1898) return "E"  ;
    if (arc_index == 1915) return "H"  ;
    if (arc_index == 1933) return "H"  ;
    if (arc_index == 1946) return "H"  ;
    if (arc_index == 1958) return "H"  ;
    if (arc_index == 1959) return "W"  ;
    if (arc_index == 1980) return "W"  ;
    if (arc_index == 1981) return "W"  ;
    if (arc_index == 1982) return "W"  ;
    if (arc_index == 1983) return "W"  ;
    if (arc_index == 1984) return "W"  ;
    if (arc_index == 1985) return "E"  ;
    if (arc_index == 1986) return "E"  ;
    if (arc_index == 1987) return "W"  ;
    if (arc_index == 1988) return "E"  ;
    if (arc_index == 1989) return "E"  ;
    if (arc_index == 1990) return "E"  ;
    if (arc_index == 1991) return "E"  ;
    if (arc_index == 1992) return "E"  ;
    if (arc_index == 1993) return "W"  ;
    if (arc_index == 1994) return "W"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 1996) return "E"  ;
    if (arc_index == 1997) return "E"  ;
    if (arc_index == 1998) return "E"  ;
    if (arc_index == 1999) return "E"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2001) return "E"  ;
    if (arc_index == 2013) return "H"  ;
    if (arc_index == 2023) return "E"  ;
    if (arc_index == 2057) return "E"  ;
    if (arc_index == 2058) return "H"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2148) return "W"  ;
    if (arc_index == 2149) return "W"  ;
    if (arc_index == 2154) return "W"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2223) return "E"  ;
    if (arc_index == 2257) return "H"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2434) return "H"  ;
    if (arc_index == 2457) return "H"  ;
    if (arc_index == 2465) return "E"  ;
    if (arc_index == 2467) return "E"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2471) return "E"  ;
    if (arc_index == 2476) return "E"  ;
    if (arc_index == 2481) return "E"  ;
    if (arc_index == 2482) return "E"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2497) return "W"  ;
    if (arc_index == 2508) return "E"  ;
    if (arc_index == 2510) return "E"  ;
    if (arc_index == 2518) return "H"  ;
    if (arc_index == 2532) return "W"  ;
    if (arc_index == 2542) return "W"  ;
    if (arc_index == 2547) return "W"  ;
    if (arc_index == 2554) return "E"  ;
    if (arc_index == 2564) return "E"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2627) return "H"  ;
    if (arc_index == 2691) return "H"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2728) return "W"  ;
    if (arc_index == 2736) return "E"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2743) return "H"  ;
    if (arc_index == 2750) return "H"  ;
    if (arc_index == 2757) return "E"  ;
    if (arc_index == 2774) return "E"  ;
    if (arc_index == 2778) return "E"  ;
    if (arc_index == 2781) return "E"  ;
    if (arc_index == 2783) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2785) return "E"  ;
    if (arc_index == 2789) return "E"  ;
    if (arc_index == 2793) return "E"  ;
    if (arc_index == 2794) return "E"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2805) return "E"  ;
    if (arc_index == 2807) return "E"  ;
    if (arc_index == 2810) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2827) return "W"  ;
    if (arc_index == 2832) return "H"  ;
    if (arc_index == 2845) return "E"  ;
    if (arc_index == 2846) return "H"  ;
    if (arc_index == 2847) return "H"  ;
    if (arc_index == 2855) return "H"  ;
    if (arc_index == 2862) return "E"  ;
    if (arc_index == 2888) return "W"  ;
    if (arc_index == 2890) return "W"  ;
    if (arc_index == 2918) return "W"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 2)) begin 
    if (arc_index == 40) return "W"  ;
    if (arc_index == 73) return "H"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 226) return "H"  ;
    if (arc_index == 407) return "W"  ;
    if (arc_index == 411) return "W"  ;
    if (arc_index == 417) return "W"  ;
    if (arc_index == 662) return "W"  ;
    if (arc_index == 681) return "W"  ;
    if (arc_index == 859) return "W"  ;
    if (arc_index == 875) return "H"  ;
    if (arc_index == 934) return "E"  ;
    if (arc_index == 936) return "E"  ;
    if (arc_index == 990) return "W"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1014) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1019) return "E"  ;
    if (arc_index == 1023) return "E"  ;
    if (arc_index == 1030) return "H"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1163) return "H"  ;
    if (arc_index == 1171) return "H"  ;
    if (arc_index == 1258) return "H"  ;
    if (arc_index == 1289) return "W"  ;
    if (arc_index == 1384) return "H"  ;
    if (arc_index == 1495) return "H"  ;
    if (arc_index == 1526) return "E"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1565) return "H"  ;
    if (arc_index == 1740) return "H"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1937) return "H"  ;
    if (arc_index == 1980) return "H"  ;
    if (arc_index == 2002) return "H"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2004) return "E"  ;
    if (arc_index == 2005) return "E"  ;
    if (arc_index == 2006) return "E"  ;
    if (arc_index == 2007) return "E"  ;
    if (arc_index == 2008) return "E"  ;
    if (arc_index == 2009) return "W"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2011) return "E"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2013) return "E"  ;
    if (arc_index == 2014) return "E"  ;
    if (arc_index == 2015) return "E"  ;
    if (arc_index == 2016) return "E"  ;
    if (arc_index == 2017) return "E"  ;
    if (arc_index == 2018) return "E"  ;
    if (arc_index == 2019) return "E"  ;
    if (arc_index == 2020) return "E"  ;
    if (arc_index == 2021) return "E"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2023) return "E"  ;
    if (arc_index == 2035) return "H"  ;
    if (arc_index == 2080) return "H"  ;
    if (arc_index == 2230) return "E"  ;
    if (arc_index == 2279) return "H"  ;
    if (arc_index == 2456) return "H"  ;
    if (arc_index == 2540) return "H"  ;
    if (arc_index == 2649) return "H"  ;
    if (arc_index == 2765) return "H"  ;
    if (arc_index == 2854) return "H"  ;
    if (arc_index == 2868) return "H"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 3)) begin 
    if (arc_index == 26) return "H"  ;
    if (arc_index == 95) return "H"  ;
    if (arc_index == 247) return "H"  ;
    if (arc_index == 248) return "H"  ;
    if (arc_index == 256) return "W"  ;
    if (arc_index == 340) return "W"  ;
    if (arc_index == 450) return "W"  ;
    if (arc_index == 472) return "W"  ;
    if (arc_index == 486) return "E"  ;
    if (arc_index == 493) return "E"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 664) return "E"  ;
    if (arc_index == 675) return "E"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 751) return "W"  ;
    if (arc_index == 753) return "W"  ;
    if (arc_index == 766) return "W"  ;
    if (arc_index == 775) return "E"  ;
    if (arc_index == 785) return "E"  ;
    if (arc_index == 848) return "W"  ;
    if (arc_index == 889) return "E"  ;
    if (arc_index == 897) return "H"  ;
    if (arc_index == 909) return "H"  ;
    if (arc_index == 950) return "E"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 1052) return "H"  ;
    if (arc_index == 1120) return "W"  ;
    if (arc_index == 1185) return "H"  ;
    if (arc_index == 1193) return "H"  ;
    if (arc_index == 1202) return "E"  ;
    if (arc_index == 1280) return "H"  ;
    if (arc_index == 1308) return "H"  ;
    if (arc_index == 1389) return "H"  ;
    if (arc_index == 1400) return "H"  ;
    if (arc_index == 1406) return "H"  ;
    if (arc_index == 1424) return "W"  ;
    if (arc_index == 1454) return "W"  ;
    if (arc_index == 1476) return "W"  ;
    if (arc_index == 1517) return "H"  ;
    if (arc_index == 1587) return "H"  ;
    if (arc_index == 1600) return "E"  ;
    if (arc_index == 1622) return "W"  ;
    if (arc_index == 1629) return "E"  ;
    if (arc_index == 1706) return "W"  ;
    if (arc_index == 1709) return "W"  ;
    if (arc_index == 1712) return "W"  ;
    if (arc_index == 1738) return "E"  ;
    if (arc_index == 1745) return "E"  ;
    if (arc_index == 1751) return "E"  ;
    if (arc_index == 1755) return "E"  ;
    if (arc_index == 1757) return "E"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1762) return "H"  ;
    if (arc_index == 1771) return "W"  ;
    if (arc_index == 1816) return "W"  ;
    if (arc_index == 1838) return "E"  ;
    if (arc_index == 1840) return "E"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1941) return "W"  ;
    if (arc_index == 1959) return "H"  ;
    if (arc_index == 2002) return "H"  ;
    if (arc_index == 2007) return "H"  ;
    if (arc_index == 2024) return "H"  ;
    if (arc_index == 2025) return "E"  ;
    if (arc_index == 2026) return "E"  ;
    if (arc_index == 2027) return "E"  ;
    if (arc_index == 2028) return "E"  ;
    if (arc_index == 2029) return "W"  ;
    if (arc_index == 2030) return "W"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2032) return "E"  ;
    if (arc_index == 2033) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2035) return "E"  ;
    if (arc_index == 2036) return "E"  ;
    if (arc_index == 2037) return "E"  ;
    if (arc_index == 2038) return "E"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2040) return "E"  ;
    if (arc_index == 2041) return "E"  ;
    if (arc_index == 2042) return "E"  ;
    if (arc_index == 2043) return "E"  ;
    if (arc_index == 2044) return "E"  ;
    if (arc_index == 2045) return "E"  ;
    if (arc_index == 2057) return "H"  ;
    if (arc_index == 2102) return "H"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2291) return "W"  ;
    if (arc_index == 2297) return "W"  ;
    if (arc_index == 2301) return "H"  ;
    if (arc_index == 2305) return "W"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2478) return "H"  ;
    if (arc_index == 2501) return "W"  ;
    if (arc_index == 2562) return "H"  ;
    if (arc_index == 2564) return "E"  ;
    if (arc_index == 2565) return "E"  ;
    if (arc_index == 2576) return "E"  ;
    if (arc_index == 2597) return "E"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2604) return "W"  ;
    if (arc_index == 2671) return "H"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2702) return "E"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2728) return "E"  ;
    if (arc_index == 2731) return "E"  ;
    if (arc_index == 2732) return "E"  ;
    if (arc_index == 2736) return "E"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2742) return "E"  ;
    if (arc_index == 2744) return "E"  ;
    if (arc_index == 2749) return "E"  ;
    if (arc_index == 2772) return "E"  ;
    if (arc_index == 2780) return "E"  ;
    if (arc_index == 2787) return "H"  ;
    if (arc_index == 2788) return "H"  ;
    if (arc_index == 2792) return "H"  ;
    if (arc_index == 2840) return "H"  ;
    if (arc_index == 2841) return "E"  ;
    if (arc_index == 2842) return "E"  ;
    if (arc_index == 2854) return "E"  ;
    if (arc_index == 2856) return "E"  ;
    if (arc_index == 2864) return "E"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2873) return "E"  ;
    if (arc_index == 2876) return "H"  ;
    if (arc_index == 2890) return "H"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 4)) begin 
    if (arc_index == 25) return "W"  ;
    if (arc_index == 26) return "W"  ;
    if (arc_index == 28) return "W"  ;
    if (arc_index == 34) return "W"  ;
    if (arc_index == 49) return "W"  ;
    if (arc_index == 50) return "W"  ;
    if (arc_index == 51) return "W"  ;
    if (arc_index == 58) return "W"  ;
    if (arc_index == 63) return "W"  ;
    if (arc_index == 65) return "W"  ;
    if (arc_index == 70) return "W"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 78) return "E"  ;
    if (arc_index == 81) return "E"  ;
    if (arc_index == 84) return "E"  ;
    if (arc_index == 86) return "E"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 117) return "H"  ;
    if (arc_index == 123) return "H"  ;
    if (arc_index == 136) return "H"  ;
    if (arc_index == 142) return "H"  ;
    if (arc_index == 185) return "H"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 270) return "H"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 284) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 362) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 410) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 456) return "E"  ;
    if (arc_index == 463) return "E"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 468) return "E"  ;
    if (arc_index == 469) return "E"  ;
    if (arc_index == 474) return "E"  ;
    if (arc_index == 476) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 481) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 540) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 656) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 726) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 752) return "W"  ;
    if (arc_index == 785) return "W"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 837) return "W"  ;
    if (arc_index == 862) return "W"  ;
    if (arc_index == 888) return "W"  ;
    if (arc_index == 890) return "E"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 895) return "E"  ;
    if (arc_index == 896) return "E"  ;
    if (arc_index == 904) return "E"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 911) return "E"  ;
    if (arc_index == 917) return "E"  ;
    if (arc_index == 919) return "H"  ;
    if (arc_index == 920) return "E"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 972) return "E"  ;
    if (arc_index == 980) return "W"  ;
    if (arc_index == 987) return "W"  ;
    if (arc_index == 988) return "W"  ;
    if (arc_index == 996) return "W"  ;
    if (arc_index == 1005) return "W"  ;
    if (arc_index == 1008) return "W"  ;
    if (arc_index == 1009) return "W"  ;
    if (arc_index == 1017) return "E"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1044) return "E"  ;
    if (arc_index == 1047) return "E"  ;
    if (arc_index == 1068) return "W"  ;
    if (arc_index == 1074) return "H"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1109) return "W"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1169) return "W"  ;
    if (arc_index == 1185) return "W"  ;
    if (arc_index == 1197) return "W"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1207) return "H"  ;
    if (arc_index == 1215) return "H"  ;
    if (arc_index == 1230) return "H"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1296) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1302) return "H"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1328) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1390) return "W"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1428) return "H"  ;
    if (arc_index == 1438) return "W"  ;
    if (arc_index == 1440) return "W"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1539) return "H"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1605) return "E"  ;
    if (arc_index == 1609) return "H"  ;
    if (arc_index == 1611) return "H"  ;
    if (arc_index == 1627) return "H"  ;
    if (arc_index == 1640) return "H"  ;
    if (arc_index == 1648) return "H"  ;
    if (arc_index == 1660) return "H"  ;
    if (arc_index == 1674) return "H"  ;
    if (arc_index == 1676) return "W"  ;
    if (arc_index == 1683) return "W"  ;
    if (arc_index == 1690) return "W"  ;
    if (arc_index == 1697) return "W"  ;
    if (arc_index == 1698) return "W"  ;
    if (arc_index == 1731) return "W"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1776) return "E"  ;
    if (arc_index == 1784) return "H"  ;
    if (arc_index == 1785) return "W"  ;
    if (arc_index == 1789) return "W"  ;
    if (arc_index == 1834) return "W"  ;
    if (arc_index == 1843) return "W"  ;
    if (arc_index == 1856) return "W"  ;
    if (arc_index == 1857) return "W"  ;
    if (arc_index == 1865) return "W"  ;
    if (arc_index == 1883) return "W"  ;
    if (arc_index == 1894) return "W"  ;
    if (arc_index == 1899) return "W"  ;
    if (arc_index == 1913) return "W"  ;
    if (arc_index == 1923) return "W"  ;
    if (arc_index == 1938) return "W"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1949) return "E"  ;
    if (arc_index == 1960) return "W"  ;
    if (arc_index == 1972) return "W"  ;
    if (arc_index == 1980) return "W"  ;
    if (arc_index == 1981) return "H"  ;
    if (arc_index == 1983) return "H"  ;
    if (arc_index == 1998) return "H"  ;
    if (arc_index == 2006) return "H"  ;
    if (arc_index == 2012) return "H"  ;
    if (arc_index == 2024) return "H"  ;
    if (arc_index == 2039) return "H"  ;
    if (arc_index == 2046) return "E"  ;
    if (arc_index == 2047) return "E"  ;
    if (arc_index == 2048) return "E"  ;
    if (arc_index == 2049) return "E"  ;
    if (arc_index == 2050) return "E"  ;
    if (arc_index == 2051) return "E"  ;
    if (arc_index == 2052) return "W"  ;
    if (arc_index == 2053) return "W"  ;
    if (arc_index == 2054) return "W"  ;
    if (arc_index == 2055) return "W"  ;
    if (arc_index == 2056) return "W"  ;
    if (arc_index == 2057) return "W"  ;
    if (arc_index == 2058) return "W"  ;
    if (arc_index == 2059) return "W"  ;
    if (arc_index == 2060) return "W"  ;
    if (arc_index == 2061) return "W"  ;
    if (arc_index == 2062) return "W"  ;
    if (arc_index == 2063) return "E"  ;
    if (arc_index == 2064) return "E"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2066) return "W"  ;
    if (arc_index == 2067) return "W"  ;
    if (arc_index == 2079) return "H"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2091) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2116) return "W"  ;
    if (arc_index == 2124) return "H"  ;
    if (arc_index == 2131) return "H"  ;
    if (arc_index == 2138) return "H"  ;
    if (arc_index == 2144) return "H"  ;
    if (arc_index == 2148) return "H"  ;
    if (arc_index == 2149) return "H"  ;
    if (arc_index == 2152) return "H"  ;
    if (arc_index == 2154) return "H"  ;
    if (arc_index == 2160) return "H"  ;
    if (arc_index == 2172) return "E"  ;
    if (arc_index == 2222) return "E"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2235) return "E"  ;
    if (arc_index == 2236) return "E"  ;
    if (arc_index == 2237) return "E"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2243) return "E"  ;
    if (arc_index == 2248) return "W"  ;
    if (arc_index == 2255) return "W"  ;
    if (arc_index == 2261) return "W"  ;
    if (arc_index == 2323) return "H"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2416) return "W"  ;
    if (arc_index == 2424) return "W"  ;
    if (arc_index == 2429) return "W"  ;
    if (arc_index == 2432) return "E"  ;
    if (arc_index == 2445) return "E"  ;
    if (arc_index == 2451) return "E"  ;
    if (arc_index == 2457) return "E"  ;
    if (arc_index == 2458) return "E"  ;
    if (arc_index == 2475) return "E"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2500) return "H"  ;
    if (arc_index == 2510) return "H"  ;
    if (arc_index == 2518) return "H"  ;
    if (arc_index == 2519) return "H"  ;
    if (arc_index == 2535) return "W"  ;
    if (arc_index == 2541) return "W"  ;
    if (arc_index == 2549) return "W"  ;
    if (arc_index == 2566) return "E"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2584) return "H"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2664) return "W"  ;
    if (arc_index == 2669) return "E"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2686) return "E"  ;
    if (arc_index == 2693) return "H"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2752) return "E"  ;
    if (arc_index == 2774) return "E"  ;
    if (arc_index == 2781) return "E"  ;
    if (arc_index == 2785) return "E"  ;
    if (arc_index == 2789) return "E"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2809) return "H"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2883) return "E"  ;
    if (arc_index == 2884) return "E"  ;
    if (arc_index == 2885) return "E"  ;
    if (arc_index == 2887) return "W"  ;
    if (arc_index == 2891) return "E"  ;
    if (arc_index == 2896) return "E"  ;
    if (arc_index == 2897) return "E"  ;
    if (arc_index == 2898) return "H"  ;
    if (arc_index == 2912) return "H"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 10)) begin 
    if (arc_index == 8) return "H"  ;
    if (arc_index == 139) return "H"  ;
    if (arc_index == 146) return "H"  ;
    if (arc_index == 283) return "H"  ;
    if (arc_index == 289) return "H"  ;
    if (arc_index == 291) return "H"  ;
    if (arc_index == 292) return "H"  ;
    if (arc_index == 370) return "H"  ;
    if (arc_index == 427) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 614) return "W"  ;
    if (arc_index == 615) return "W"  ;
    if (arc_index == 685) return "W"  ;
    if (arc_index == 723) return "W"  ;
    if (arc_index == 740) return "W"  ;
    if (arc_index == 818) return "W"  ;
    if (arc_index == 941) return "H"  ;
    if (arc_index == 1037) return "H"  ;
    if (arc_index == 1053) return "H"  ;
    if (arc_index == 1057) return "H"  ;
    if (arc_index == 1096) return "H"  ;
    if (arc_index == 1100) return "H"  ;
    if (arc_index == 1122) return "H"  ;
    if (arc_index == 1124) return "H"  ;
    if (arc_index == 1127) return "H"  ;
    if (arc_index == 1128) return "H"  ;
    if (arc_index == 1130) return "H"  ;
    if (arc_index == 1132) return "H"  ;
    if (arc_index == 1133) return "H"  ;
    if (arc_index == 1134) return "H"  ;
    if (arc_index == 1136) return "H"  ;
    if (arc_index == 1138) return "H"  ;
    if (arc_index == 1140) return "H"  ;
    if (arc_index == 1141) return "H"  ;
    if (arc_index == 1142) return "H"  ;
    if (arc_index == 1143) return "H"  ;
    if (arc_index == 1155) return "H"  ;
    if (arc_index == 1229) return "H"  ;
    if (arc_index == 1237) return "H"  ;
    if (arc_index == 1241) return "H"  ;
    if (arc_index == 1249) return "H"  ;
    if (arc_index == 1324) return "H"  ;
    if (arc_index == 1399) return "H"  ;
    if (arc_index == 1450) return "H"  ;
    if (arc_index == 1540) return "H"  ;
    if (arc_index == 1561) return "H"  ;
    if (arc_index == 1567) return "H"  ;
    if (arc_index == 1570) return "H"  ;
    if (arc_index == 1577) return "H"  ;
    if (arc_index == 1579) return "E"  ;
    if (arc_index == 1580) return "E"  ;
    if (arc_index == 1583) return "E"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1631) return "H"  ;
    if (arc_index == 1660) return "H"  ;
    if (arc_index == 1668) return "H"  ;
    if (arc_index == 1769) return "H"  ;
    if (arc_index == 1806) return "H"  ;
    if (arc_index == 1839) return "H"  ;
    if (arc_index == 2003) return "H"  ;
    if (arc_index == 2046) return "H"  ;
    if (arc_index == 2068) return "H"  ;
    if (arc_index == 2069) return "W"  ;
    if (arc_index == 2070) return "W"  ;
    if (arc_index == 2071) return "W"  ;
    if (arc_index == 2072) return "W"  ;
    if (arc_index == 2073) return "W"  ;
    if (arc_index == 2074) return "W"  ;
    if (arc_index == 2075) return "W"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2077) return "W"  ;
    if (arc_index == 2078) return "W"  ;
    if (arc_index == 2079) return "W"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2081) return "W"  ;
    if (arc_index == 2082) return "W"  ;
    if (arc_index == 2083) return "W"  ;
    if (arc_index == 2084) return "W"  ;
    if (arc_index == 2085) return "W"  ;
    if (arc_index == 2086) return "W"  ;
    if (arc_index == 2087) return "W"  ;
    if (arc_index == 2088) return "W"  ;
    if (arc_index == 2089) return "W"  ;
    if (arc_index == 2100) return "W"  ;
    if (arc_index == 2101) return "H"  ;
    if (arc_index == 2146) return "H"  ;
    if (arc_index == 2178) return "H"  ;
    if (arc_index == 2184) return "H"  ;
    if (arc_index == 2197) return "W"  ;
    if (arc_index == 2208) return "W"  ;
    if (arc_index == 2211) return "W"  ;
    if (arc_index == 2345) return "H"  ;
    if (arc_index == 2382) return "W"  ;
    if (arc_index == 2396) return "W"  ;
    if (arc_index == 2414) return "W"  ;
    if (arc_index == 2522) return "H"  ;
    if (arc_index == 2559) return "H"  ;
    if (arc_index == 2595) return "H"  ;
    if (arc_index == 2606) return "H"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2712) return "W"  ;
    if (arc_index == 2715) return "H"  ;
    if (arc_index == 2831) return "H"  ;
    if (arc_index == 2920) return "H"  ;
    if (arc_index == 2921) return "H"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 8)) begin 
    if (arc_index == 16) return "H"  ;
    if (arc_index == 30) return "H"  ;
    if (arc_index == 161) return "H"  ;
    if (arc_index == 314) return "H"  ;
    if (arc_index == 528) return "W"  ;
    if (arc_index == 551) return "E"  ;
    if (arc_index == 552) return "E"  ;
    if (arc_index == 556) return "E"  ;
    if (arc_index == 558) return "E"  ;
    if (arc_index == 563) return "E"  ;
    if (arc_index == 566) return "E"  ;
    if (arc_index == 568) return "E"  ;
    if (arc_index == 628) return "W"  ;
    if (arc_index == 788) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 963) return "H"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1118) return "H"  ;
    if (arc_index == 1251) return "H"  ;
    if (arc_index == 1259) return "H"  ;
    if (arc_index == 1343) return "W"  ;
    if (arc_index == 1346) return "H"  ;
    if (arc_index == 1426) return "H"  ;
    if (arc_index == 1472) return "H"  ;
    if (arc_index == 1498) return "E"  ;
    if (arc_index == 1547) return "W"  ;
    if (arc_index == 1583) return "H"  ;
    if (arc_index == 1653) return "H"  ;
    if (arc_index == 1695) return "E"  ;
    if (arc_index == 1701) return "E"  ;
    if (arc_index == 1708) return "E"  ;
    if (arc_index == 1738) return "E"  ;
    if (arc_index == 1760) return "E"  ;
    if (arc_index == 1761) return "W"  ;
    if (arc_index == 1762) return "W"  ;
    if (arc_index == 1763) return "W"  ;
    if (arc_index == 1764) return "W"  ;
    if (arc_index == 1767) return "W"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1771) return "W"  ;
    if (arc_index == 1772) return "W"  ;
    if (arc_index == 1773) return "W"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1778) return "W"  ;
    if (arc_index == 1781) return "W"  ;
    if (arc_index == 1793) return "E"  ;
    if (arc_index == 1828) return "H"  ;
    if (arc_index == 1838) return "E"  ;
    if (arc_index == 2025) return "H"  ;
    if (arc_index == 2037) return "E"  ;
    if (arc_index == 2068) return "H"  ;
    if (arc_index == 2090) return "H"  ;
    if (arc_index == 2091) return "H"  ;
    if (arc_index == 2092) return "H"  ;
    if (arc_index == 2093) return "H"  ;
    if (arc_index == 2094) return "W"  ;
    if (arc_index == 2095) return "W"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2097) return "W"  ;
    if (arc_index == 2098) return "W"  ;
    if (arc_index == 2099) return "W"  ;
    if (arc_index == 2100) return "W"  ;
    if (arc_index == 2101) return "E"  ;
    if (arc_index == 2102) return "W"  ;
    if (arc_index == 2103) return "W"  ;
    if (arc_index == 2104) return "W"  ;
    if (arc_index == 2105) return "E"  ;
    if (arc_index == 2106) return "E"  ;
    if (arc_index == 2107) return "E"  ;
    if (arc_index == 2108) return "E"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2110) return "W"  ;
    if (arc_index == 2111) return "E"  ;
    if (arc_index == 2123) return "H"  ;
    if (arc_index == 2168) return "H"  ;
    if (arc_index == 2214) return "E"  ;
    if (arc_index == 2298) return "E"  ;
    if (arc_index == 2349) return "W"  ;
    if (arc_index == 2367) return "H"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2544) return "H"  ;
    if (arc_index == 2572) return "H"  ;
    if (arc_index == 2628) return "H"  ;
    if (arc_index == 2737) return "H"  ;
    if (arc_index == 2853) return "H"  ;
    if (arc_index == 2916) return "W"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 5)) begin 
    if (arc_index == 0) return "W"  ;
    if (arc_index == 30) return "W"  ;
    if (arc_index == 38) return "H"  ;
    if (arc_index == 52) return "H"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 72) return "E"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 78) return "E"  ;
    if (arc_index == 81) return "E"  ;
    if (arc_index == 84) return "E"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 98) return "E"  ;
    if (arc_index == 101) return "E"  ;
    if (arc_index == 116) return "E"  ;
    if (arc_index == 123) return "W"  ;
    if (arc_index == 125) return "E"  ;
    if (arc_index == 130) return "E"  ;
    if (arc_index == 159) return "E"  ;
    if (arc_index == 183) return "H"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 210) return "W"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 270) return "W"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 284) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 336) return "H"  ;
    if (arc_index == 367) return "H"  ;
    if (arc_index == 373) return "H"  ;
    if (arc_index == 386) return "H"  ;
    if (arc_index == 399) return "H"  ;
    if (arc_index == 403) return "E"  ;
    if (arc_index == 412) return "E"  ;
    if (arc_index == 414) return "E"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 455) return "E"  ;
    if (arc_index == 463) return "E"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 468) return "E"  ;
    if (arc_index == 469) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 481) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 502) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 525) return "E"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 656) return "W"  ;
    if (arc_index == 663) return "W"  ;
    if (arc_index == 686) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 691) return "W"  ;
    if (arc_index == 726) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 757) return "W"  ;
    if (arc_index == 759) return "W"  ;
    if (arc_index == 769) return "W"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 829) return "E"  ;
    if (arc_index == 837) return "W"  ;
    if (arc_index == 862) return "W"  ;
    if (arc_index == 876) return "W"  ;
    if (arc_index == 879) return "W"  ;
    if (arc_index == 890) return "E"  ;
    if (arc_index == 904) return "E"  ;
    if (arc_index == 905) return "E"  ;
    if (arc_index == 911) return "E"  ;
    if (arc_index == 917) return "E"  ;
    if (arc_index == 920) return "E"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 971) return "E"  ;
    if (arc_index == 974) return "E"  ;
    if (arc_index == 980) return "W"  ;
    if (arc_index == 985) return "H"  ;
    if (arc_index == 988) return "W"  ;
    if (arc_index == 991) return "E"  ;
    if (arc_index == 1017) return "E"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1053) return "W"  ;
    if (arc_index == 1074) return "W"  ;
    if (arc_index == 1092) return "E"  ;
    if (arc_index == 1096) return "E"  ;
    if (arc_index == 1109) return "W"  ;
    if (arc_index == 1140) return "H"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1185) return "W"  ;
    if (arc_index == 1195) return "E"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1273) return "H"  ;
    if (arc_index == 1279) return "H"  ;
    if (arc_index == 1281) return "H"  ;
    if (arc_index == 1296) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1302) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1328) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1368) return "H"  ;
    if (arc_index == 1385) return "H"  ;
    if (arc_index == 1393) return "H"  ;
    if (arc_index == 1408) return "H"  ;
    if (arc_index == 1422) return "H"  ;
    if (arc_index == 1430) return "H"  ;
    if (arc_index == 1432) return "H"  ;
    if (arc_index == 1441) return "H"  ;
    if (arc_index == 1463) return "H"  ;
    if (arc_index == 1470) return "H"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1494) return "H"  ;
    if (arc_index == 1498) return "H"  ;
    if (arc_index == 1514) return "H"  ;
    if (arc_index == 1520) return "H"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1605) return "H"  ;
    if (arc_index == 1607) return "E"  ;
    if (arc_index == 1608) return "E"  ;
    if (arc_index == 1615) return "E"  ;
    if (arc_index == 1621) return "E"  ;
    if (arc_index == 1626) return "E"  ;
    if (arc_index == 1635) return "E"  ;
    if (arc_index == 1674) return "W"  ;
    if (arc_index == 1675) return "H"  ;
    if (arc_index == 1676) return "W"  ;
    if (arc_index == 1683) return "W"  ;
    if (arc_index == 1690) return "W"  ;
    if (arc_index == 1698) return "W"  ;
    if (arc_index == 1707) return "W"  ;
    if (arc_index == 1710) return "W"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1773) return "E"  ;
    if (arc_index == 1775) return "E"  ;
    if (arc_index == 1785) return "W"  ;
    if (arc_index == 1789) return "W"  ;
    if (arc_index == 1802) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1850) return "H"  ;
    if (arc_index == 1855) return "H"  ;
    if (arc_index == 1856) return "W"  ;
    if (arc_index == 1864) return "W"  ;
    if (arc_index == 1865) return "W"  ;
    if (arc_index == 1870) return "W"  ;
    if (arc_index == 1881) return "W"  ;
    if (arc_index == 1883) return "W"  ;
    if (arc_index == 1900) return "W"  ;
    if (arc_index == 1902) return "W"  ;
    if (arc_index == 1909) return "W"  ;
    if (arc_index == 1913) return "W"  ;
    if (arc_index == 1916) return "E"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1949) return "E"  ;
    if (arc_index == 1960) return "W"  ;
    if (arc_index == 1969) return "W"  ;
    if (arc_index == 1970) return "W"  ;
    if (arc_index == 1972) return "W"  ;
    if (arc_index == 1973) return "W"  ;
    if (arc_index == 2032) return "E"  ;
    if (arc_index == 2046) return "E"  ;
    if (arc_index == 2047) return "H"  ;
    if (arc_index == 2063) return "E"  ;
    if (arc_index == 2079) return "W"  ;
    if (arc_index == 2090) return "H"  ;
    if (arc_index == 2091) return "W"  ;
    if (arc_index == 2112) return "W"  ;
    if (arc_index == 2113) return "W"  ;
    if (arc_index == 2114) return "E"  ;
    if (arc_index == 2115) return "E"  ;
    if (arc_index == 2116) return "W"  ;
    if (arc_index == 2117) return "W"  ;
    if (arc_index == 2118) return "W"  ;
    if (arc_index == 2119) return "W"  ;
    if (arc_index == 2120) return "W"  ;
    if (arc_index == 2121) return "W"  ;
    if (arc_index == 2122) return "W"  ;
    if (arc_index == 2123) return "W"  ;
    if (arc_index == 2124) return "W"  ;
    if (arc_index == 2125) return "W"  ;
    if (arc_index == 2126) return "E"  ;
    if (arc_index == 2127) return "E"  ;
    if (arc_index == 2128) return "E"  ;
    if (arc_index == 2129) return "E"  ;
    if (arc_index == 2130) return "E"  ;
    if (arc_index == 2131) return "W"  ;
    if (arc_index == 2132) return "W"  ;
    if (arc_index == 2133) return "W"  ;
    if (arc_index == 2145) return "H"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2169) return "E"  ;
    if (arc_index == 2172) return "E"  ;
    if (arc_index == 2188) return "E"  ;
    if (arc_index == 2190) return "H"  ;
    if (arc_index == 2191) return "H"  ;
    if (arc_index == 2202) return "H"  ;
    if (arc_index == 2222) return "E"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2235) return "E"  ;
    if (arc_index == 2237) return "E"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2248) return "W"  ;
    if (arc_index == 2255) return "W"  ;
    if (arc_index == 2261) return "W"  ;
    if (arc_index == 2276) return "W"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2323) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2389) return "H"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2416) return "W"  ;
    if (arc_index == 2430) return "W"  ;
    if (arc_index == 2432) return "E"  ;
    if (arc_index == 2449) return "E"  ;
    if (arc_index == 2451) return "E"  ;
    if (arc_index == 2491) return "E"  ;
    if (arc_index == 2493) return "E"  ;
    if (arc_index == 2498) return "E"  ;
    if (arc_index == 2500) return "W"  ;
    if (arc_index == 2505) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2533) return "E"  ;
    if (arc_index == 2534) return "E"  ;
    if (arc_index == 2549) return "W"  ;
    if (arc_index == 2551) return "W"  ;
    if (arc_index == 2566) return "H"  ;
    if (arc_index == 2610) return "H"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2650) return "H"  ;
    if (arc_index == 2655) return "H"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2669) return "E"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2698) return "E"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2736) return "E"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2752) return "E"  ;
    if (arc_index == 2759) return "H"  ;
    if (arc_index == 2764) return "H"  ;
    if (arc_index == 2767) return "H"  ;
    if (arc_index == 2771) return "H"  ;
    if (arc_index == 2815) return "H"  ;
    if (arc_index == 2841) return "H"  ;
    if (arc_index == 2875) return "H"  ;
    if (arc_index == 2884) return "E"  ;
    if (arc_index == 2891) return "E"  ;
    if (arc_index == 2912) return "W"  ;
    if (arc_index == 2919) return "W"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 4)) begin 
    if (arc_index == 27) return "W"  ;
    if (arc_index == 36) return "W"  ;
    if (arc_index == 40) return "W"  ;
    if (arc_index == 45) return "E"  ;
    if (arc_index == 48) return "E"  ;
    if (arc_index == 54) return "E"  ;
    if (arc_index == 60) return "H"  ;
    if (arc_index == 66) return "E"  ;
    if (arc_index == 67) return "E"  ;
    if (arc_index == 74) return "H"  ;
    if (arc_index == 93) return "W"  ;
    if (arc_index == 96) return "W"  ;
    if (arc_index == 99) return "W"  ;
    if (arc_index == 102) return "W"  ;
    if (arc_index == 110) return "W"  ;
    if (arc_index == 112) return "W"  ;
    if (arc_index == 115) return "W"  ;
    if (arc_index == 120) return "W"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 135) return "W"  ;
    if (arc_index == 136) return "W"  ;
    if (arc_index == 138) return "W"  ;
    if (arc_index == 142) return "W"  ;
    if (arc_index == 145) return "W"  ;
    if (arc_index == 148) return "W"  ;
    if (arc_index == 149) return "E"  ;
    if (arc_index == 152) return "E"  ;
    if (arc_index == 163) return "E"  ;
    if (arc_index == 165) return "E"  ;
    if (arc_index == 173) return "E"  ;
    if (arc_index == 180) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 205) return "H"  ;
    if (arc_index == 210) return "H"  ;
    if (arc_index == 279) return "H"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 345) return "W"  ;
    if (arc_index == 352) return "W"  ;
    if (arc_index == 357) return "W"  ;
    if (arc_index == 358) return "H"  ;
    if (arc_index == 360) return "W"  ;
    if (arc_index == 374) return "E"  ;
    if (arc_index == 376) return "E"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 382) return "E"  ;
    if (arc_index == 385) return "E"  ;
    if (arc_index == 387) return "E"  ;
    if (arc_index == 393) return "E"  ;
    if (arc_index == 397) return "W"  ;
    if (arc_index == 405) return "W"  ;
    if (arc_index == 410) return "W"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 451) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 641) return "W"  ;
    if (arc_index == 644) return "W"  ;
    if (arc_index == 645) return "W"  ;
    if (arc_index == 651) return "W"  ;
    if (arc_index == 663) return "W"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 669) return "E"  ;
    if (arc_index == 752) return "E"  ;
    if (arc_index == 779) return "E"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 795) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 895) return "W"  ;
    if (arc_index == 915) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 940) return "E"  ;
    if (arc_index == 941) return "E"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 1001) return "E"  ;
    if (arc_index == 1007) return "H"  ;
    if (arc_index == 1014) return "H"  ;
    if (arc_index == 1019) return "H"  ;
    if (arc_index == 1020) return "H"  ;
    if (arc_index == 1033) return "H"  ;
    if (arc_index == 1041) return "H"  ;
    if (arc_index == 1131) return "H"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1162) return "H"  ;
    if (arc_index == 1204) return "H"  ;
    if (arc_index == 1240) return "W"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1267) return "W"  ;
    if (arc_index == 1282) return "W"  ;
    if (arc_index == 1289) return "W"  ;
    if (arc_index == 1295) return "H"  ;
    if (arc_index == 1303) return "H"  ;
    if (arc_index == 1378) return "W"  ;
    if (arc_index == 1390) return "H"  ;
    if (arc_index == 1423) return "H"  ;
    if (arc_index == 1439) return "W"  ;
    if (arc_index == 1470) return "W"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1516) return "H"  ;
    if (arc_index == 1529) return "E"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1603) return "W"  ;
    if (arc_index == 1611) return "W"  ;
    if (arc_index == 1627) return "H"  ;
    if (arc_index == 1677) return "W"  ;
    if (arc_index == 1687) return "W"  ;
    if (arc_index == 1697) return "H"  ;
    if (arc_index == 1698) return "H"  ;
    if (arc_index == 1723) return "E"  ;
    if (arc_index == 1724) return "E"  ;
    if (arc_index == 1764) return "W"  ;
    if (arc_index == 1775) return "W"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1824) return "W"  ;
    if (arc_index == 1856) return "W"  ;
    if (arc_index == 1872) return "H"  ;
    if (arc_index == 1878) return "W"  ;
    if (arc_index == 1890) return "W"  ;
    if (arc_index == 1931) return "W"  ;
    if (arc_index == 1935) return "W"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1980) return "E"  ;
    if (arc_index == 2004) return "E"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2069) return "H"  ;
    if (arc_index == 2071) return "W"  ;
    if (arc_index == 2074) return "W"  ;
    if (arc_index == 2112) return "H"  ;
    if (arc_index == 2134) return "W"  ;
    if (arc_index == 2135) return "E"  ;
    if (arc_index == 2136) return "E"  ;
    if (arc_index == 2137) return "E"  ;
    if (arc_index == 2138) return "E"  ;
    if (arc_index == 2139) return "E"  ;
    if (arc_index == 2140) return "W"  ;
    if (arc_index == 2141) return "W"  ;
    if (arc_index == 2142) return "E"  ;
    if (arc_index == 2143) return "E"  ;
    if (arc_index == 2144) return "E"  ;
    if (arc_index == 2145) return "E"  ;
    if (arc_index == 2146) return "E"  ;
    if (arc_index == 2147) return "E"  ;
    if (arc_index == 2148) return "E"  ;
    if (arc_index == 2149) return "E"  ;
    if (arc_index == 2150) return "E"  ;
    if (arc_index == 2151) return "E"  ;
    if (arc_index == 2152) return "E"  ;
    if (arc_index == 2153) return "E"  ;
    if (arc_index == 2154) return "E"  ;
    if (arc_index == 2155) return "E"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2167) return "H"  ;
    if (arc_index == 2175) return "E"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2212) return "H"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2227) return "W"  ;
    if (arc_index == 2246) return "W"  ;
    if (arc_index == 2279) return "W"  ;
    if (arc_index == 2411) return "H"  ;
    if (arc_index == 2420) return "H"  ;
    if (arc_index == 2437) return "E"  ;
    if (arc_index == 2445) return "E"  ;
    if (arc_index == 2451) return "E"  ;
    if (arc_index == 2452) return "E"  ;
    if (arc_index == 2457) return "E"  ;
    if (arc_index == 2458) return "E"  ;
    if (arc_index == 2460) return "E"  ;
    if (arc_index == 2463) return "E"  ;
    if (arc_index == 2475) return "E"  ;
    if (arc_index == 2483) return "E"  ;
    if (arc_index == 2510) return "E"  ;
    if (arc_index == 2512) return "E"  ;
    if (arc_index == 2517) return "E"  ;
    if (arc_index == 2518) return "E"  ;
    if (arc_index == 2519) return "E"  ;
    if (arc_index == 2521) return "E"  ;
    if (arc_index == 2522) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2524) return "E"  ;
    if (arc_index == 2525) return "E"  ;
    if (arc_index == 2528) return "E"  ;
    if (arc_index == 2529) return "E"  ;
    if (arc_index == 2551) return "E"  ;
    if (arc_index == 2588) return "H"  ;
    if (arc_index == 2592) return "E"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2672) return "H"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2719) return "E"  ;
    if (arc_index == 2733) return "E"  ;
    if (arc_index == 2781) return "H"  ;
    if (arc_index == 2796) return "H"  ;
    if (arc_index == 2812) return "H"  ;
    if (arc_index == 2885) return "E"  ;
    if (arc_index == 2896) return "E"  ;
    if (arc_index == 2897) return "H"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 3)) begin 
    if (arc_index == 1) return "W"  ;
    if (arc_index == 3) return "W"  ;
    if (arc_index == 18) return "W"  ;
    if (arc_index == 35) return "W"  ;
    if (arc_index == 41) return "W"  ;
    if (arc_index == 44) return "W"  ;
    if (arc_index == 47) return "W"  ;
    if (arc_index == 59) return "W"  ;
    if (arc_index == 61) return "W"  ;
    if (arc_index == 66) return "W"  ;
    if (arc_index == 68) return "E"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 72) return "E"  ;
    if (arc_index == 74) return "E"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 77) return "E"  ;
    if (arc_index == 78) return "E"  ;
    if (arc_index == 81) return "E"  ;
    if (arc_index == 82) return "H"  ;
    if (arc_index == 84) return "H"  ;
    if (arc_index == 86) return "H"  ;
    if (arc_index == 87) return "E"  ;
    if (arc_index == 96) return "H"  ;
    if (arc_index == 106) return "W"  ;
    if (arc_index == 107) return "W"  ;
    if (arc_index == 138) return "W"  ;
    if (arc_index == 148) return "W"  ;
    if (arc_index == 152) return "W"  ;
    if (arc_index == 159) return "W"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 222) return "W"  ;
    if (arc_index == 227) return "H"  ;
    if (arc_index == 238) return "H"  ;
    if (arc_index == 246) return "H"  ;
    if (arc_index == 268) return "H"  ;
    if (arc_index == 343) return "W"  ;
    if (arc_index == 349) return "W"  ;
    if (arc_index == 380) return "H"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 397) return "E"  ;
    if (arc_index == 404) return "E"  ;
    if (arc_index == 405) return "E"  ;
    if (arc_index == 419) return "W"  ;
    if (arc_index == 445) return "E"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 448) return "E"  ;
    if (arc_index == 458) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 461) return "E"  ;
    if (arc_index == 466) return "E"  ;
    if (arc_index == 483) return "E"  ;
    if (arc_index == 490) return "E"  ;
    if (arc_index == 496) return "E"  ;
    if (arc_index == 497) return "E"  ;
    if (arc_index == 498) return "E"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 530) return "W"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 553) return "W"  ;
    if (arc_index == 562) return "W"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 573) return "W"  ;
    if (arc_index == 579) return "W"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 582) return "E"  ;
    if (arc_index == 591) return "E"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 664) return "W"  ;
    if (arc_index == 668) return "W"  ;
    if (arc_index == 674) return "E"  ;
    if (arc_index == 675) return "E"  ;
    if (arc_index == 676) return "E"  ;
    if (arc_index == 678) return "E"  ;
    if (arc_index == 693) return "E"  ;
    if (arc_index == 703) return "E"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 750) return "W"  ;
    if (arc_index == 792) return "W"  ;
    if (arc_index == 810) return "W"  ;
    if (arc_index == 811) return "W"  ;
    if (arc_index == 812) return "E"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 903) return "E"  ;
    if (arc_index == 910) return "E"  ;
    if (arc_index == 923) return "E"  ;
    if (arc_index == 928) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 946) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 962) return "E"  ;
    if (arc_index == 994) return "E"  ;
    if (arc_index == 995) return "E"  ;
    if (arc_index == 1000) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1010) return "W"  ;
    if (arc_index == 1016) return "W"  ;
    if (arc_index == 1025) return "W"  ;
    if (arc_index == 1029) return "H"  ;
    if (arc_index == 1032) return "H"  ;
    if (arc_index == 1068) return "H"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1184) return "H"  ;
    if (arc_index == 1195) return "E"  ;
    if (arc_index == 1196) return "E"  ;
    if (arc_index == 1292) return "W"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1317) return "H"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1325) return "H"  ;
    if (arc_index == 1330) return "H"  ;
    if (arc_index == 1336) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1366) return "W"  ;
    if (arc_index == 1383) return "W"  ;
    if (arc_index == 1412) return "H"  ;
    if (arc_index == 1437) return "W"  ;
    if (arc_index == 1444) return "W"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1499) return "W"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1538) return "H"  ;
    if (arc_index == 1539) return "H"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1637) return "E"  ;
    if (arc_index == 1649) return "H"  ;
    if (arc_index == 1657) return "H"  ;
    if (arc_index == 1658) return "H"  ;
    if (arc_index == 1659) return "W"  ;
    if (arc_index == 1669) return "W"  ;
    if (arc_index == 1676) return "W"  ;
    if (arc_index == 1719) return "H"  ;
    if (arc_index == 1724) return "H"  ;
    if (arc_index == 1753) return "H"  ;
    if (arc_index == 1789) return "W"  ;
    if (arc_index == 1839) return "W"  ;
    if (arc_index == 1842) return "W"  ;
    if (arc_index == 1857) return "W"  ;
    if (arc_index == 1865) return "W"  ;
    if (arc_index == 1871) return "W"  ;
    if (arc_index == 1894) return "H"  ;
    if (arc_index == 1913) return "H"  ;
    if (arc_index == 1929) return "E"  ;
    if (arc_index == 1931) return "E"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 1972) return "W"  ;
    if (arc_index == 1987) return "W"  ;
    if (arc_index == 2001) return "W"  ;
    if (arc_index == 2006) return "E"  ;
    if (arc_index == 2013) return "E"  ;
    if (arc_index == 2023) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2040) return "W"  ;
    if (arc_index == 2054) return "W"  ;
    if (arc_index == 2067) return "W"  ;
    if (arc_index == 2091) return "H"  ;
    if (arc_index == 2134) return "H"  ;
    if (arc_index == 2153) return "W"  ;
    if (arc_index == 2155) return "W"  ;
    if (arc_index == 2156) return "E"  ;
    if (arc_index == 2157) return "E"  ;
    if (arc_index == 2158) return "E"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2161) return "W"  ;
    if (arc_index == 2162) return "W"  ;
    if (arc_index == 2163) return "E"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2165) return "W"  ;
    if (arc_index == 2166) return "W"  ;
    if (arc_index == 2167) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2169) return "E"  ;
    if (arc_index == 2170) return "E"  ;
    if (arc_index == 2171) return "E"  ;
    if (arc_index == 2172) return "E"  ;
    if (arc_index == 2173) return "W"  ;
    if (arc_index == 2174) return "E"  ;
    if (arc_index == 2175) return "E"  ;
    if (arc_index == 2176) return "E"  ;
    if (arc_index == 2177) return "E"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2189) return "H"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2226) return "E"  ;
    if (arc_index == 2227) return "E"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2234) return "H"  ;
    if (arc_index == 2275) return "W"  ;
    if (arc_index == 2281) return "W"  ;
    if (arc_index == 2283) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2421) return "W"  ;
    if (arc_index == 2422) return "W"  ;
    if (arc_index == 2423) return "W"  ;
    if (arc_index == 2424) return "E"  ;
    if (arc_index == 2429) return "E"  ;
    if (arc_index == 2432) return "E"  ;
    if (arc_index == 2433) return "H"  ;
    if (arc_index == 2434) return "H"  ;
    if (arc_index == 2438) return "W"  ;
    if (arc_index == 2442) return "W"  ;
    if (arc_index == 2450) return "W"  ;
    if (arc_index == 2460) return "W"  ;
    if (arc_index == 2483) return "W"  ;
    if (arc_index == 2486) return "W"  ;
    if (arc_index == 2508) return "W"  ;
    if (arc_index == 2516) return "W"  ;
    if (arc_index == 2535) return "W"  ;
    if (arc_index == 2540) return "W"  ;
    if (arc_index == 2580) return "E"  ;
    if (arc_index == 2610) return "H"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2694) return "H"  ;
    if (arc_index == 2697) return "H"  ;
    if (arc_index == 2704) return "E"  ;
    if (arc_index == 2723) return "E"  ;
    if (arc_index == 2755) return "E"  ;
    if (arc_index == 2789) return "E"  ;
    if (arc_index == 2793) return "W"  ;
    if (arc_index == 2796) return "W"  ;
    if (arc_index == 2803) return "H"  ;
    if (arc_index == 2812) return "H"  ;
    if (arc_index == 2842) return "H"  ;
    if (arc_index == 2854) return "H"  ;
    if (arc_index == 2887) return "H"  ;
    if (arc_index == 2919) return "H"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 10)) begin 
    if (arc_index == 15) return "H"  ;
    if (arc_index == 57) return "E"  ;
    if (arc_index == 104) return "H"  ;
    if (arc_index == 118) return "H"  ;
    if (arc_index == 177) return "W"  ;
    if (arc_index == 179) return "W"  ;
    if (arc_index == 183) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 191) return "W"  ;
    if (arc_index == 196) return "W"  ;
    if (arc_index == 197) return "W"  ;
    if (arc_index == 203) return "W"  ;
    if (arc_index == 209) return "W"  ;
    if (arc_index == 234) return "E"  ;
    if (arc_index == 249) return "H"  ;
    if (arc_index == 254) return "H"  ;
    if (arc_index == 287) return "W"  ;
    if (arc_index == 289) return "W"  ;
    if (arc_index == 290) return "W"  ;
    if (arc_index == 291) return "W"  ;
    if (arc_index == 292) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 298) return "W"  ;
    if (arc_index == 303) return "W"  ;
    if (arc_index == 304) return "W"  ;
    if (arc_index == 370) return "W"  ;
    if (arc_index == 402) return "H"  ;
    if (arc_index == 543) return "E"  ;
    if (arc_index == 544) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 614) return "E"  ;
    if (arc_index == 615) return "E"  ;
    if (arc_index == 616) return "W"  ;
    if (arc_index == 620) return "W"  ;
    if (arc_index == 630) return "W"  ;
    if (arc_index == 646) return "E"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 714) return "E"  ;
    if (arc_index == 723) return "E"  ;
    if (arc_index == 740) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 818) return "E"  ;
    if (arc_index == 823) return "E"  ;
    if (arc_index == 871) return "E"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 1037) return "E"  ;
    if (arc_index == 1051) return "H"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1053) return "W"  ;
    if (arc_index == 1054) return "W"  ;
    if (arc_index == 1067) return "W"  ;
    if (arc_index == 1112) return "W"  ;
    if (arc_index == 1122) return "W"  ;
    if (arc_index == 1128) return "W"  ;
    if (arc_index == 1132) return "W"  ;
    if (arc_index == 1133) return "W"  ;
    if (arc_index == 1134) return "W"  ;
    if (arc_index == 1138) return "W"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1155) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1206) return "H"  ;
    if (arc_index == 1241) return "H"  ;
    if (arc_index == 1249) return "H"  ;
    if (arc_index == 1324) return "H"  ;
    if (arc_index == 1326) return "H"  ;
    if (arc_index == 1339) return "H"  ;
    if (arc_index == 1342) return "W"  ;
    if (arc_index == 1347) return "H"  ;
    if (arc_index == 1399) return "H"  ;
    if (arc_index == 1434) return "H"  ;
    if (arc_index == 1446) return "H"  ;
    if (arc_index == 1450) return "H"  ;
    if (arc_index == 1488) return "E"  ;
    if (arc_index == 1560) return "H"  ;
    if (arc_index == 1561) return "H"  ;
    if (arc_index == 1570) return "H"  ;
    if (arc_index == 1577) return "H"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1671) return "H"  ;
    if (arc_index == 1681) return "E"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1741) return "H"  ;
    if (arc_index == 1769) return "H"  ;
    if (arc_index == 1806) return "H"  ;
    if (arc_index == 1809) return "E"  ;
    if (arc_index == 1867) return "E"  ;
    if (arc_index == 1875) return "E"  ;
    if (arc_index == 1916) return "H"  ;
    if (arc_index == 1962) return "E"  ;
    if (arc_index == 1975) return "E"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2068) return "W"  ;
    if (arc_index == 2070) return "W"  ;
    if (arc_index == 2073) return "E"  ;
    if (arc_index == 2075) return "E"  ;
    if (arc_index == 2078) return "E"  ;
    if (arc_index == 2081) return "E"  ;
    if (arc_index == 2083) return "E"  ;
    if (arc_index == 2085) return "E"  ;
    if (arc_index == 2088) return "E"  ;
    if (arc_index == 2089) return "E"  ;
    if (arc_index == 2100) return "E"  ;
    if (arc_index == 2101) return "E"  ;
    if (arc_index == 2113) return "H"  ;
    if (arc_index == 2156) return "H"  ;
    if (arc_index == 2178) return "H"  ;
    if (arc_index == 2179) return "W"  ;
    if (arc_index == 2180) return "W"  ;
    if (arc_index == 2181) return "W"  ;
    if (arc_index == 2182) return "W"  ;
    if (arc_index == 2183) return "W"  ;
    if (arc_index == 2184) return "W"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2186) return "W"  ;
    if (arc_index == 2187) return "W"  ;
    if (arc_index == 2188) return "W"  ;
    if (arc_index == 2189) return "W"  ;
    if (arc_index == 2190) return "W"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2193) return "W"  ;
    if (arc_index == 2194) return "W"  ;
    if (arc_index == 2195) return "W"  ;
    if (arc_index == 2196) return "W"  ;
    if (arc_index == 2197) return "W"  ;
    if (arc_index == 2198) return "W"  ;
    if (arc_index == 2199) return "E"  ;
    if (arc_index == 2208) return "E"  ;
    if (arc_index == 2211) return "H"  ;
    if (arc_index == 2256) return "H"  ;
    if (arc_index == 2269) return "E"  ;
    if (arc_index == 2271) return "E"  ;
    if (arc_index == 2311) return "E"  ;
    if (arc_index == 2345) return "E"  ;
    if (arc_index == 2358) return "E"  ;
    if (arc_index == 2377) return "W"  ;
    if (arc_index == 2382) return "W"  ;
    if (arc_index == 2444) return "E"  ;
    if (arc_index == 2455) return "H"  ;
    if (arc_index == 2484) return "H"  ;
    if (arc_index == 2606) return "H"  ;
    if (arc_index == 2621) return "H"  ;
    if (arc_index == 2632) return "H"  ;
    if (arc_index == 2638) return "W"  ;
    if (arc_index == 2639) return "W"  ;
    if (arc_index == 2643) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2708) return "W"  ;
    if (arc_index == 2709) return "W"  ;
    if (arc_index == 2710) return "W"  ;
    if (arc_index == 2712) return "W"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2714) return "W"  ;
    if (arc_index == 2716) return "H"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2719) return "W"  ;
    if (arc_index == 2720) return "W"  ;
    if (arc_index == 2721) return "W"  ;
    if (arc_index == 2722) return "W"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2725) return "W"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2825) return "H"  ;
    if (arc_index == 2831) return "H"  ;
    if (arc_index == 2920) return "H"  ;
    if (arc_index == 2921) return "H"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 8)) begin 
    if (arc_index == 37) return "H"  ;
    if (arc_index == 126) return "H"  ;
    if (arc_index == 139) return "E"  ;
    if (arc_index == 140) return "H"  ;
    if (arc_index == 146) return "E"  ;
    if (arc_index == 150) return "E"  ;
    if (arc_index == 219) return "E"  ;
    if (arc_index == 240) return "E"  ;
    if (arc_index == 252) return "E"  ;
    if (arc_index == 271) return "H"  ;
    if (arc_index == 361) return "H"  ;
    if (arc_index == 364) return "H"  ;
    if (arc_index == 370) return "E"  ;
    if (arc_index == 416) return "E"  ;
    if (arc_index == 423) return "E"  ;
    if (arc_index == 424) return "H"  ;
    if (arc_index == 425) return "E"  ;
    if (arc_index == 427) return "E"  ;
    if (arc_index == 432) return "E"  ;
    if (arc_index == 435) return "E"  ;
    if (arc_index == 459) return "E"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 467) return "E"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 704) return "E"  ;
    if (arc_index == 726) return "E"  ;
    if (arc_index == 729) return "E"  ;
    if (arc_index == 730) return "E"  ;
    if (arc_index == 733) return "E"  ;
    if (arc_index == 734) return "E"  ;
    if (arc_index == 735) return "W"  ;
    if (arc_index == 736) return "W"  ;
    if (arc_index == 737) return "W"  ;
    if (arc_index == 739) return "W"  ;
    if (arc_index == 740) return "W"  ;
    if (arc_index == 741) return "W"  ;
    if (arc_index == 742) return "W"  ;
    if (arc_index == 743) return "W"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 747) return "W"  ;
    if (arc_index == 759) return "W"  ;
    if (arc_index == 825) return "W"  ;
    if (arc_index == 860) return "E"  ;
    if (arc_index == 867) return "E"  ;
    if (arc_index == 1012) return "E"  ;
    if (arc_index == 1041) return "W"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1045) return "W"  ;
    if (arc_index == 1046) return "W"  ;
    if (arc_index == 1073) return "H"  ;
    if (arc_index == 1123) return "W"  ;
    if (arc_index == 1129) return "W"  ;
    if (arc_index == 1131) return "W"  ;
    if (arc_index == 1135) return "W"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1139) return "W"  ;
    if (arc_index == 1228) return "H"  ;
    if (arc_index == 1264) return "H"  ;
    if (arc_index == 1270) return "W"  ;
    if (arc_index == 1276) return "E"  ;
    if (arc_index == 1299) return "W"  ;
    if (arc_index == 1307) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1312) return "W"  ;
    if (arc_index == 1314) return "W"  ;
    if (arc_index == 1315) return "W"  ;
    if (arc_index == 1317) return "W"  ;
    if (arc_index == 1318) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1361) return "H"  ;
    if (arc_index == 1369) return "H"  ;
    if (arc_index == 1376) return "E"  ;
    if (arc_index == 1456) return "H"  ;
    if (arc_index == 1489) return "H"  ;
    if (arc_index == 1497) return "H"  ;
    if (arc_index == 1501) return "H"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1574) return "W"  ;
    if (arc_index == 1582) return "H"  ;
    if (arc_index == 1693) return "H"  ;
    if (arc_index == 1763) return "H"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1876) return "E"  ;
    if (arc_index == 1885) return "E"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 1938) return "H"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1988) return "E"  ;
    if (arc_index == 2017) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2061) return "E"  ;
    if (arc_index == 2080) return "W"  ;
    if (arc_index == 2086) return "W"  ;
    if (arc_index == 2119) return "E"  ;
    if (arc_index == 2135) return "H"  ;
    if (arc_index == 2150) return "E"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2178) return "H"  ;
    if (arc_index == 2180) return "W"  ;
    if (arc_index == 2200) return "W"  ;
    if (arc_index == 2201) return "W"  ;
    if (arc_index == 2202) return "W"  ;
    if (arc_index == 2203) return "E"  ;
    if (arc_index == 2204) return "W"  ;
    if (arc_index == 2205) return "W"  ;
    if (arc_index == 2206) return "W"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2208) return "W"  ;
    if (arc_index == 2209) return "W"  ;
    if (arc_index == 2210) return "W"  ;
    if (arc_index == 2211) return "E"  ;
    if (arc_index == 2212) return "W"  ;
    if (arc_index == 2213) return "W"  ;
    if (arc_index == 2214) return "W"  ;
    if (arc_index == 2215) return "W"  ;
    if (arc_index == 2216) return "W"  ;
    if (arc_index == 2217) return "W"  ;
    if (arc_index == 2218) return "W"  ;
    if (arc_index == 2219) return "W"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2233) return "H"  ;
    if (arc_index == 2278) return "H"  ;
    if (arc_index == 2314) return "W"  ;
    if (arc_index == 2361) return "W"  ;
    if (arc_index == 2377) return "W"  ;
    if (arc_index == 2428) return "W"  ;
    if (arc_index == 2448) return "E"  ;
    if (arc_index == 2455) return "E"  ;
    if (arc_index == 2462) return "E"  ;
    if (arc_index == 2477) return "H"  ;
    if (arc_index == 2525) return "H"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2621) return "E"  ;
    if (arc_index == 2640) return "E"  ;
    if (arc_index == 2646) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2654) return "H"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2680) return "W"  ;
    if (arc_index == 2726) return "W"  ;
    if (arc_index == 2738) return "H"  ;
    if (arc_index == 2821) return "H"  ;
    if (arc_index == 2847) return "H"  ;
    if (arc_index == 2908) return "H"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 1)) begin 
    if (arc_index == 13) return "W"  ;
    if (arc_index == 59) return "H"  ;
    if (arc_index == 69) return "H"  ;
    if (arc_index == 145) return "H"  ;
    if (arc_index == 148) return "H"  ;
    if (arc_index == 162) return "H"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 274) return "W"  ;
    if (arc_index == 293) return "H"  ;
    if (arc_index == 384) return "H"  ;
    if (arc_index == 388) return "W"  ;
    if (arc_index == 389) return "W"  ;
    if (arc_index == 440) return "E"  ;
    if (arc_index == 441) return "E"  ;
    if (arc_index == 446) return "H"  ;
    if (arc_index == 449) return "H"  ;
    if (arc_index == 450) return "H"  ;
    if (arc_index == 460) return "H"  ;
    if (arc_index == 462) return "H"  ;
    if (arc_index == 473) return "H"  ;
    if (arc_index == 484) return "H"  ;
    if (arc_index == 495) return "E"  ;
    if (arc_index == 501) return "E"  ;
    if (arc_index == 513) return "E"  ;
    if (arc_index == 514) return "E"  ;
    if (arc_index == 517) return "E"  ;
    if (arc_index == 518) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 582) return "E"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 641) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 773) return "W"  ;
    if (arc_index == 774) return "W"  ;
    if (arc_index == 800) return "W"  ;
    if (arc_index == 809) return "W"  ;
    if (arc_index == 886) return "W"  ;
    if (arc_index == 894) return "W"  ;
    if (arc_index == 924) return "W"  ;
    if (arc_index == 948) return "W"  ;
    if (arc_index == 957) return "W"  ;
    if (arc_index == 979) return "W"  ;
    if (arc_index == 1013) return "W"  ;
    if (arc_index == 1017) return "E"  ;
    if (arc_index == 1018) return "E"  ;
    if (arc_index == 1024) return "E"  ;
    if (arc_index == 1087) return "E"  ;
    if (arc_index == 1090) return "E"  ;
    if (arc_index == 1095) return "H"  ;
    if (arc_index == 1145) return "H"  ;
    if (arc_index == 1213) return "E"  ;
    if (arc_index == 1223) return "E"  ;
    if (arc_index == 1224) return "E"  ;
    if (arc_index == 1225) return "E"  ;
    if (arc_index == 1250) return "H"  ;
    if (arc_index == 1318) return "H"  ;
    if (arc_index == 1372) return "H"  ;
    if (arc_index == 1383) return "H"  ;
    if (arc_index == 1391) return "H"  ;
    if (arc_index == 1478) return "H"  ;
    if (arc_index == 1499) return "H"  ;
    if (arc_index == 1527) return "E"  ;
    if (arc_index == 1532) return "E"  ;
    if (arc_index == 1590) return "E"  ;
    if (arc_index == 1604) return "H"  ;
    if (arc_index == 1634) return "H"  ;
    if (arc_index == 1664) return "H"  ;
    if (arc_index == 1690) return "W"  ;
    if (arc_index == 1715) return "H"  ;
    if (arc_index == 1748) return "H"  ;
    if (arc_index == 1785) return "H"  ;
    if (arc_index == 1823) return "W"  ;
    if (arc_index == 1830) return "W"  ;
    if (arc_index == 1831) return "W"  ;
    if (arc_index == 1937) return "W"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1942) return "E"  ;
    if (arc_index == 1945) return "E"  ;
    if (arc_index == 1950) return "E"  ;
    if (arc_index == 1951) return "E"  ;
    if (arc_index == 1956) return "E"  ;
    if (arc_index == 1960) return "H"  ;
    if (arc_index == 2014) return "H"  ;
    if (arc_index == 2021) return "H"  ;
    if (arc_index == 2116) return "H"  ;
    if (arc_index == 2155) return "W"  ;
    if (arc_index == 2157) return "H"  ;
    if (arc_index == 2176) return "H"  ;
    if (arc_index == 2200) return "H"  ;
    if (arc_index == 2213) return "H"  ;
    if (arc_index == 2221) return "H"  ;
    if (arc_index == 2222) return "E"  ;
    if (arc_index == 2223) return "E"  ;
    if (arc_index == 2224) return "E"  ;
    if (arc_index == 2225) return "W"  ;
    if (arc_index == 2226) return "W"  ;
    if (arc_index == 2227) return "E"  ;
    if (arc_index == 2228) return "E"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2230) return "E"  ;
    if (arc_index == 2231) return "W"  ;
    if (arc_index == 2232) return "W"  ;
    if (arc_index == 2233) return "E"  ;
    if (arc_index == 2234) return "E"  ;
    if (arc_index == 2235) return "E"  ;
    if (arc_index == 2236) return "E"  ;
    if (arc_index == 2237) return "E"  ;
    if (arc_index == 2238) return "E"  ;
    if (arc_index == 2239) return "E"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2241) return "E"  ;
    if (arc_index == 2242) return "E"  ;
    if (arc_index == 2243) return "E"  ;
    if (arc_index == 2255) return "H"  ;
    if (arc_index == 2300) return "H"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2423) return "W"  ;
    if (arc_index == 2450) return "W"  ;
    if (arc_index == 2499) return "H"  ;
    if (arc_index == 2552) return "H"  ;
    if (arc_index == 2556) return "H"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2576) return "E"  ;
    if (arc_index == 2582) return "E"  ;
    if (arc_index == 2583) return "E"  ;
    if (arc_index == 2585) return "E"  ;
    if (arc_index == 2593) return "E"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2662) return "E"  ;
    if (arc_index == 2664) return "E"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2669) return "E"  ;
    if (arc_index == 2670) return "E"  ;
    if (arc_index == 2672) return "E"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2676) return "H"  ;
    if (arc_index == 2677) return "E"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2682) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2730) return "E"  ;
    if (arc_index == 2747) return "E"  ;
    if (arc_index == 2748) return "E"  ;
    if (arc_index == 2760) return "H"  ;
    if (arc_index == 2796) return "E"  ;
    if (arc_index == 2811) return "E"  ;
    if (arc_index == 2851) return "E"  ;
    if (arc_index == 2859) return "E"  ;
    if (arc_index == 2863) return "E"  ;
    if (arc_index == 2869) return "H"  ;
    if (arc_index == 2874) return "H"  ;
    if (arc_index == 2879) return "H"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 6)) begin 
    if (arc_index == 1) return "H"  ;
    if (arc_index == 3) return "H"  ;
    if (arc_index == 19) return "H"  ;
    if (arc_index == 20) return "H"  ;
    if (arc_index == 33) return "H"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 64) return "E"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 81) return "H"  ;
    if (arc_index == 84) return "H"  ;
    if (arc_index == 98) return "W"  ;
    if (arc_index == 101) return "W"  ;
    if (arc_index == 113) return "W"  ;
    if (arc_index == 125) return "W"  ;
    if (arc_index == 128) return "W"  ;
    if (arc_index == 132) return "E"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 170) return "H"  ;
    if (arc_index == 173) return "H"  ;
    if (arc_index == 183) return "W"  ;
    if (arc_index == 184) return "H"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 205) return "W"  ;
    if (arc_index == 210) return "W"  ;
    if (arc_index == 265) return "W"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 270) return "W"  ;
    if (arc_index == 284) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 308) return "W"  ;
    if (arc_index == 315) return "H"  ;
    if (arc_index == 327) return "H"  ;
    if (arc_index == 332) return "H"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 338) return "E"  ;
    if (arc_index == 340) return "E"  ;
    if (arc_index == 342) return "E"  ;
    if (arc_index == 344) return "E"  ;
    if (arc_index == 347) return "E"  ;
    if (arc_index == 356) return "E"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 403) return "W"  ;
    if (arc_index == 426) return "W"  ;
    if (arc_index == 436) return "W"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 463) return "E"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 468) return "H"  ;
    if (arc_index == 469) return "E"  ;
    if (arc_index == 477) return "E"  ;
    if (arc_index == 481) return "E"  ;
    if (arc_index == 489) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 535) return "E"  ;
    if (arc_index == 564) return "E"  ;
    if (arc_index == 607) return "E"  ;
    if (arc_index == 629) return "E"  ;
    if (arc_index == 642) return "E"  ;
    if (arc_index == 647) return "E"  ;
    if (arc_index == 649) return "E"  ;
    if (arc_index == 653) return "E"  ;
    if (arc_index == 654) return "E"  ;
    if (arc_index == 655) return "E"  ;
    if (arc_index == 656) return "W"  ;
    if (arc_index == 667) return "W"  ;
    if (arc_index == 677) return "E"  ;
    if (arc_index == 691) return "W"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 784) return "W"  ;
    if (arc_index == 791) return "W"  ;
    if (arc_index == 792) return "E"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 836) return "W"  ;
    if (arc_index == 839) return "W"  ;
    if (arc_index == 850) return "W"  ;
    if (arc_index == 851) return "W"  ;
    if (arc_index == 863) return "W"  ;
    if (arc_index == 866) return "W"  ;
    if (arc_index == 869) return "W"  ;
    if (arc_index == 876) return "W"  ;
    if (arc_index == 890) return "W"  ;
    if (arc_index == 898) return "W"  ;
    if (arc_index == 905) return "W"  ;
    if (arc_index == 911) return "E"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 928) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 991) return "E"  ;
    if (arc_index == 997) return "E"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1053) return "W"  ;
    if (arc_index == 1059) return "W"  ;
    if (arc_index == 1074) return "W"  ;
    if (arc_index == 1085) return "W"  ;
    if (arc_index == 1092) return "W"  ;
    if (arc_index == 1093) return "W"  ;
    if (arc_index == 1100) return "W"  ;
    if (arc_index == 1101) return "W"  ;
    if (arc_index == 1102) return "W"  ;
    if (arc_index == 1107) return "W"  ;
    if (arc_index == 1109) return "W"  ;
    if (arc_index == 1112) return "E"  ;
    if (arc_index == 1114) return "E"  ;
    if (arc_index == 1115) return "E"  ;
    if (arc_index == 1117) return "H"  ;
    if (arc_index == 1124) return "H"  ;
    if (arc_index == 1140) return "W"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1170) return "W"  ;
    if (arc_index == 1174) return "W"  ;
    if (arc_index == 1178) return "W"  ;
    if (arc_index == 1185) return "W"  ;
    if (arc_index == 1186) return "E"  ;
    if (arc_index == 1187) return "E"  ;
    if (arc_index == 1195) return "E"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1272) return "H"  ;
    if (arc_index == 1273) return "W"  ;
    if (arc_index == 1275) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1302) return "W"  ;
    if (arc_index == 1325) return "W"  ;
    if (arc_index == 1327) return "W"  ;
    if (arc_index == 1328) return "W"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1377) return "W"  ;
    if (arc_index == 1396) return "W"  ;
    if (arc_index == 1397) return "W"  ;
    if (arc_index == 1401) return "W"  ;
    if (arc_index == 1405) return "H"  ;
    if (arc_index == 1413) return "H"  ;
    if (arc_index == 1415) return "H"  ;
    if (arc_index == 1449) return "H"  ;
    if (arc_index == 1456) return "H"  ;
    if (arc_index == 1462) return "H"  ;
    if (arc_index == 1470) return "W"  ;
    if (arc_index == 1471) return "W"  ;
    if (arc_index == 1480) return "W"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1490) return "W"  ;
    if (arc_index == 1500) return "H"  ;
    if (arc_index == 1507) return "H"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1607) return "E"  ;
    if (arc_index == 1608) return "E"  ;
    if (arc_index == 1620) return "E"  ;
    if (arc_index == 1626) return "H"  ;
    if (arc_index == 1641) return "H"  ;
    if (arc_index == 1650) return "E"  ;
    if (arc_index == 1671) return "E"  ;
    if (arc_index == 1674) return "W"  ;
    if (arc_index == 1675) return "W"  ;
    if (arc_index == 1676) return "W"  ;
    if (arc_index == 1683) return "W"  ;
    if (arc_index == 1684) return "W"  ;
    if (arc_index == 1687) return "W"  ;
    if (arc_index == 1690) return "W"  ;
    if (arc_index == 1691) return "W"  ;
    if (arc_index == 1704) return "W"  ;
    if (arc_index == 1730) return "E"  ;
    if (arc_index == 1737) return "H"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1788) return "E"  ;
    if (arc_index == 1807) return "H"  ;
    if (arc_index == 1813) return "H"  ;
    if (arc_index == 1820) return "H"  ;
    if (arc_index == 1821) return "H"  ;
    if (arc_index == 1848) return "H"  ;
    if (arc_index == 1870) return "W"  ;
    if (arc_index == 1896) return "W"  ;
    if (arc_index == 1916) return "W"  ;
    if (arc_index == 1949) return "E"  ;
    if (arc_index == 1960) return "W"  ;
    if (arc_index == 1965) return "W"  ;
    if (arc_index == 1968) return "W"  ;
    if (arc_index == 1969) return "W"  ;
    if (arc_index == 1970) return "W"  ;
    if (arc_index == 1972) return "W"  ;
    if (arc_index == 1973) return "W"  ;
    if (arc_index == 1982) return "H"  ;
    if (arc_index == 1988) return "H"  ;
    if (arc_index == 2031) return "H"  ;
    if (arc_index == 2032) return "H"  ;
    if (arc_index == 2046) return "E"  ;
    if (arc_index == 2063) return "E"  ;
    if (arc_index == 2079) return "W"  ;
    if (arc_index == 2114) return "E"  ;
    if (arc_index == 2126) return "E"  ;
    if (arc_index == 2129) return "E"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2172) return "E"  ;
    if (arc_index == 2179) return "H"  ;
    if (arc_index == 2188) return "W"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2222) return "H"  ;
    if (arc_index == 2233) return "H"  ;
    if (arc_index == 2235) return "E"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2244) return "E"  ;
    if (arc_index == 2245) return "E"  ;
    if (arc_index == 2246) return "E"  ;
    if (arc_index == 2247) return "E"  ;
    if (arc_index == 2248) return "W"  ;
    if (arc_index == 2249) return "W"  ;
    if (arc_index == 2250) return "W"  ;
    if (arc_index == 2251) return "W"  ;
    if (arc_index == 2252) return "W"  ;
    if (arc_index == 2253) return "W"  ;
    if (arc_index == 2254) return "W"  ;
    if (arc_index == 2255) return "W"  ;
    if (arc_index == 2256) return "W"  ;
    if (arc_index == 2257) return "W"  ;
    if (arc_index == 2258) return "W"  ;
    if (arc_index == 2259) return "W"  ;
    if (arc_index == 2260) return "W"  ;
    if (arc_index == 2261) return "W"  ;
    if (arc_index == 2262) return "W"  ;
    if (arc_index == 2263) return "W"  ;
    if (arc_index == 2264) return "W"  ;
    if (arc_index == 2265) return "W"  ;
    if (arc_index == 2274) return "W"  ;
    if (arc_index == 2276) return "W"  ;
    if (arc_index == 2277) return "H"  ;
    if (arc_index == 2280) return "H"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2322) return "H"  ;
    if (arc_index == 2323) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2389) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2398) return "W"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2416) return "W"  ;
    if (arc_index == 2432) return "E"  ;
    if (arc_index == 2451) return "E"  ;
    if (arc_index == 2505) return "E"  ;
    if (arc_index == 2521) return "H"  ;
    if (arc_index == 2614) return "H"  ;
    if (arc_index == 2622) return "H"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2669) return "E"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2698) return "H"  ;
    if (arc_index == 2705) return "E"  ;
    if (arc_index == 2707) return "E"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2736) return "W"  ;
    if (arc_index == 2738) return "W"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2749) return "E"  ;
    if (arc_index == 2782) return "H"  ;
    if (arc_index == 2813) return "H"  ;
    if (arc_index == 2819) return "H"  ;
    if (arc_index == 2820) return "H"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2884) return "E"  ;
    if (arc_index == 2891) return "H"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 7)) begin 
    if (arc_index == 21) return "E"  ;
    if (arc_index == 29) return "E"  ;
    if (arc_index == 43) return "E"  ;
    if (arc_index == 53) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 57) return "E"  ;
    if (arc_index == 62) return "E"  ;
    if (arc_index == 91) return "E"  ;
    if (arc_index == 92) return "E"  ;
    if (arc_index == 95) return "E"  ;
    if (arc_index == 97) return "E"  ;
    if (arc_index == 101) return "E"  ;
    if (arc_index == 103) return "H"  ;
    if (arc_index == 109) return "E"  ;
    if (arc_index == 118) return "E"  ;
    if (arc_index == 119) return "E"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 156) return "E"  ;
    if (arc_index == 165) return "W"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 176) return "W"  ;
    if (arc_index == 182) return "W"  ;
    if (arc_index == 184) return "W"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 192) return "H"  ;
    if (arc_index == 201) return "W"  ;
    if (arc_index == 206) return "H"  ;
    if (arc_index == 222) return "W"  ;
    if (arc_index == 223) return "W"  ;
    if (arc_index == 224) return "W"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 227) return "W"  ;
    if (arc_index == 238) return "W"  ;
    if (arc_index == 257) return "W"  ;
    if (arc_index == 299) return "W"  ;
    if (arc_index == 303) return "W"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 337) return "H"  ;
    if (arc_index == 339) return "E"  ;
    if (arc_index == 341) return "E"  ;
    if (arc_index == 348) return "E"  ;
    if (arc_index == 354) return "E"  ;
    if (arc_index == 359) return "E"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 402) return "E"  ;
    if (arc_index == 428) return "E"  ;
    if (arc_index == 431) return "E"  ;
    if (arc_index == 433) return "E"  ;
    if (arc_index == 438) return "E"  ;
    if (arc_index == 463) return "E"  ;
    if (arc_index == 464) return "E"  ;
    if (arc_index == 490) return "H"  ;
    if (arc_index == 496) return "H"  ;
    if (arc_index == 497) return "E"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 530) return "W"  ;
    if (arc_index == 533) return "W"  ;
    if (arc_index == 535) return "W"  ;
    if (arc_index == 540) return "W"  ;
    if (arc_index == 546) return "W"  ;
    if (arc_index == 561) return "E"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 595) return "E"  ;
    if (arc_index == 599) return "W"  ;
    if (arc_index == 604) return "W"  ;
    if (arc_index == 639) return "E"  ;
    if (arc_index == 643) return "E"  ;
    if (arc_index == 652) return "E"  ;
    if (arc_index == 660) return "E"  ;
    if (arc_index == 674) return "E"  ;
    if (arc_index == 695) return "E"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 733) return "W"  ;
    if (arc_index == 742) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 769) return "W"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 828) return "E"  ;
    if (arc_index == 839) return "E"  ;
    if (arc_index == 851) return "E"  ;
    if (arc_index == 857) return "E"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 973) return "E"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 983) return "E"  ;
    if (arc_index == 986) return "E"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1035) return "E"  ;
    if (arc_index == 1053) return "E"  ;
    if (arc_index == 1057) return "E"  ;
    if (arc_index == 1065) return "E"  ;
    if (arc_index == 1069) return "E"  ;
    if (arc_index == 1072) return "E"  ;
    if (arc_index == 1112) return "E"  ;
    if (arc_index == 1124) return "E"  ;
    if (arc_index == 1127) return "E"  ;
    if (arc_index == 1139) return "H"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1144) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1163) return "W"  ;
    if (arc_index == 1175) return "E"  ;
    if (arc_index == 1177) return "E"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1214) return "E"  ;
    if (arc_index == 1217) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1250) return "W"  ;
    if (arc_index == 1269) return "W"  ;
    if (arc_index == 1273) return "W"  ;
    if (arc_index == 1277) return "W"  ;
    if (arc_index == 1280) return "W"  ;
    if (arc_index == 1281) return "W"  ;
    if (arc_index == 1286) return "W"  ;
    if (arc_index == 1290) return "W"  ;
    if (arc_index == 1291) return "E"  ;
    if (arc_index == 1294) return "H"  ;
    if (arc_index == 1297) return "H"  ;
    if (arc_index == 1302) return "H"  ;
    if (arc_index == 1306) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1354) return "W"  ;
    if (arc_index == 1364) return "W"  ;
    if (arc_index == 1367) return "W"  ;
    if (arc_index == 1374) return "W"  ;
    if (arc_index == 1375) return "W"  ;
    if (arc_index == 1379) return "W"  ;
    if (arc_index == 1380) return "E"  ;
    if (arc_index == 1385) return "W"  ;
    if (arc_index == 1397) return "W"  ;
    if (arc_index == 1415) return "W"  ;
    if (arc_index == 1427) return "H"  ;
    if (arc_index == 1434) return "E"  ;
    if (arc_index == 1435) return "H"  ;
    if (arc_index == 1436) return "E"  ;
    if (arc_index == 1445) return "E"  ;
    if (arc_index == 1446) return "E"  ;
    if (arc_index == 1450) return "E"  ;
    if (arc_index == 1451) return "E"  ;
    if (arc_index == 1474) return "W"  ;
    if (arc_index == 1510) return "W"  ;
    if (arc_index == 1515) return "W"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1522) return "H"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1546) return "E"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1553) return "W"  ;
    if (arc_index == 1608) return "W"  ;
    if (arc_index == 1641) return "W"  ;
    if (arc_index == 1648) return "H"  ;
    if (arc_index == 1730) return "H"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1759) return "H"  ;
    if (arc_index == 1764) return "W"  ;
    if (arc_index == 1801) return "W"  ;
    if (arc_index == 1803) return "W"  ;
    if (arc_index == 1810) return "W"  ;
    if (arc_index == 1814) return "W"  ;
    if (arc_index == 1818) return "W"  ;
    if (arc_index == 1829) return "H"  ;
    if (arc_index == 1848) return "H"  ;
    if (arc_index == 1877) return "H"  ;
    if (arc_index == 1889) return "H"  ;
    if (arc_index == 1900) return "H"  ;
    if (arc_index == 1916) return "E"  ;
    if (arc_index == 1938) return "E"  ;
    if (arc_index == 1976) return "E"  ;
    if (arc_index == 2004) return "H"  ;
    if (arc_index == 2010) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2042) return "E"  ;
    if (arc_index == 2046) return "E"  ;
    if (arc_index == 2048) return "E"  ;
    if (arc_index == 2077) return "W"  ;
    if (arc_index == 2087) return "W"  ;
    if (arc_index == 2113) return "E"  ;
    if (arc_index == 2128) return "E"  ;
    if (arc_index == 2141) return "E"  ;
    if (arc_index == 2156) return "E"  ;
    if (arc_index == 2174) return "E"  ;
    if (arc_index == 2179) return "W"  ;
    if (arc_index == 2185) return "W"  ;
    if (arc_index == 2189) return "W"  ;
    if (arc_index == 2190) return "W"  ;
    if (arc_index == 2193) return "W"  ;
    if (arc_index == 2201) return "H"  ;
    if (arc_index == 2206) return "H"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2244) return "H"  ;
    if (arc_index == 2245) return "E"  ;
    if (arc_index == 2256) return "E"  ;
    if (arc_index == 2263) return "E"  ;
    if (arc_index == 2266) return "E"  ;
    if (arc_index == 2267) return "E"  ;
    if (arc_index == 2268) return "E"  ;
    if (arc_index == 2269) return "E"  ;
    if (arc_index == 2270) return "E"  ;
    if (arc_index == 2271) return "E"  ;
    if (arc_index == 2272) return "E"  ;
    if (arc_index == 2273) return "E"  ;
    if (arc_index == 2274) return "W"  ;
    if (arc_index == 2275) return "W"  ;
    if (arc_index == 2276) return "W"  ;
    if (arc_index == 2277) return "W"  ;
    if (arc_index == 2278) return "E"  ;
    if (arc_index == 2279) return "W"  ;
    if (arc_index == 2280) return "W"  ;
    if (arc_index == 2281) return "W"  ;
    if (arc_index == 2282) return "W"  ;
    if (arc_index == 2283) return "W"  ;
    if (arc_index == 2284) return "W"  ;
    if (arc_index == 2285) return "W"  ;
    if (arc_index == 2286) return "W"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2296) return "W"  ;
    if (arc_index == 2299) return "H"  ;
    if (arc_index == 2306) return "W"  ;
    if (arc_index == 2318) return "W"  ;
    if (arc_index == 2321) return "W"  ;
    if (arc_index == 2323) return "W"  ;
    if (arc_index == 2344) return "H"  ;
    if (arc_index == 2348) return "H"  ;
    if (arc_index == 2350) return "H"  ;
    if (arc_index == 2372) return "H"  ;
    if (arc_index == 2417) return "W"  ;
    if (arc_index == 2418) return "W"  ;
    if (arc_index == 2431) return "E"  ;
    if (arc_index == 2435) return "E"  ;
    if (arc_index == 2446) return "E"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2507) return "E"  ;
    if (arc_index == 2524) return "E"  ;
    if (arc_index == 2543) return "H"  ;
    if (arc_index == 2559) return "H"  ;
    if (arc_index == 2638) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2708) return "W"  ;
    if (arc_index == 2720) return "H"  ;
    if (arc_index == 2721) return "H"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2764) return "E"  ;
    if (arc_index == 2804) return "H"  ;
    if (arc_index == 2821) return "E"  ;
    if (arc_index == 2837) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2884) return "E"  ;
    if (arc_index == 2905) return "W"  ;
    if (arc_index == 2913) return "H"  ;
    if (arc_index == 2922) return "H"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 7)) begin 
    if (arc_index == 9) return "H"  ;
    if (arc_index == 16) return "E"  ;
    if (arc_index == 43) return "E"  ;
    if (arc_index == 86) return "E"  ;
    if (arc_index == 125) return "H"  ;
    if (arc_index == 164) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 214) return "H"  ;
    if (arc_index == 228) return "H"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 247) return "W"  ;
    if (arc_index == 248) return "W"  ;
    if (arc_index == 251) return "W"  ;
    if (arc_index == 256) return "W"  ;
    if (arc_index == 259) return "W"  ;
    if (arc_index == 262) return "W"  ;
    if (arc_index == 263) return "W"  ;
    if (arc_index == 281) return "W"  ;
    if (arc_index == 288) return "W"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 359) return "H"  ;
    if (arc_index == 512) return "H"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 554) return "E"  ;
    if (arc_index == 557) return "E"  ;
    if (arc_index == 561) return "E"  ;
    if (arc_index == 564) return "E"  ;
    if (arc_index == 621) return "W"  ;
    if (arc_index == 683) return "W"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 708) return "W"  ;
    if (arc_index == 712) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 719) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 722) return "W"  ;
    if (arc_index == 749) return "W"  ;
    if (arc_index == 780) return "E"  ;
    if (arc_index == 782) return "E"  ;
    if (arc_index == 827) return "E"  ;
    if (arc_index == 834) return "W"  ;
    if (arc_index == 889) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1088) return "E"  ;
    if (arc_index == 1094) return "E"  ;
    if (arc_index == 1108) return "E"  ;
    if (arc_index == 1146) return "W"  ;
    if (arc_index == 1161) return "H"  ;
    if (arc_index == 1313) return "H"  ;
    if (arc_index == 1316) return "H"  ;
    if (arc_index == 1392) return "E"  ;
    if (arc_index == 1402) return "E"  ;
    if (arc_index == 1409) return "E"  ;
    if (arc_index == 1420) return "E"  ;
    if (arc_index == 1449) return "H"  ;
    if (arc_index == 1457) return "H"  ;
    if (arc_index == 1458) return "E"  ;
    if (arc_index == 1467) return "E"  ;
    if (arc_index == 1468) return "E"  ;
    if (arc_index == 1469) return "E"  ;
    if (arc_index == 1486) return "W"  ;
    if (arc_index == 1544) return "H"  ;
    if (arc_index == 1624) return "E"  ;
    if (arc_index == 1670) return "H"  ;
    if (arc_index == 1685) return "W"  ;
    if (arc_index == 1705) return "E"  ;
    if (arc_index == 1714) return "E"  ;
    if (arc_index == 1738) return "E"  ;
    if (arc_index == 1757) return "E"  ;
    if (arc_index == 1758) return "E"  ;
    if (arc_index == 1760) return "W"  ;
    if (arc_index == 1764) return "W"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1773) return "W"  ;
    if (arc_index == 1781) return "H"  ;
    if (arc_index == 1828) return "E"  ;
    if (arc_index == 1851) return "H"  ;
    if (arc_index == 1854) return "E"  ;
    if (arc_index == 2026) return "H"  ;
    if (arc_index == 2041) return "E"  ;
    if (arc_index == 2099) return "W"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2223) return "H"  ;
    if (arc_index == 2266) return "H"  ;
    if (arc_index == 2288) return "H"  ;
    if (arc_index == 2289) return "E"  ;
    if (arc_index == 2290) return "W"  ;
    if (arc_index == 2291) return "W"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2293) return "W"  ;
    if (arc_index == 2294) return "W"  ;
    if (arc_index == 2295) return "W"  ;
    if (arc_index == 2296) return "W"  ;
    if (arc_index == 2297) return "W"  ;
    if (arc_index == 2298) return "W"  ;
    if (arc_index == 2299) return "W"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2301) return "W"  ;
    if (arc_index == 2302) return "W"  ;
    if (arc_index == 2303) return "W"  ;
    if (arc_index == 2304) return "W"  ;
    if (arc_index == 2305) return "W"  ;
    if (arc_index == 2306) return "W"  ;
    if (arc_index == 2307) return "W"  ;
    if (arc_index == 2308) return "W"  ;
    if (arc_index == 2309) return "W"  ;
    if (arc_index == 2321) return "H"  ;
    if (arc_index == 2335) return "H"  ;
    if (arc_index == 2341) return "H"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2366) return "H"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2503) return "E"  ;
    if (arc_index == 2504) return "E"  ;
    if (arc_index == 2531) return "E"  ;
    if (arc_index == 2550) return "E"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2565) return "H"  ;
    if (arc_index == 2570) return "H"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2602) return "W"  ;
    if (arc_index == 2603) return "W"  ;
    if (arc_index == 2604) return "W"  ;
    if (arc_index == 2608) return "W"  ;
    if (arc_index == 2617) return "W"  ;
    if (arc_index == 2637) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2731) return "E"  ;
    if (arc_index == 2742) return "H"  ;
    if (arc_index == 2776) return "H"  ;
    if (arc_index == 2777) return "H"  ;
    if (arc_index == 2791) return "E"  ;
    if (arc_index == 2816) return "W"  ;
    if (arc_index == 2826) return "H"  ;
    if (arc_index == 2829) return "W"  ;
    if (arc_index == 2864) return "W"  ;
    if (arc_index == 2870) return "W"  ;
    if (arc_index == 2873) return "E"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 9)) begin 
    if (arc_index == 8) return "E"  ;
    if (arc_index == 31) return "H"  ;
    if (arc_index == 62) return "E"  ;
    if (arc_index == 104) return "E"  ;
    if (arc_index == 111) return "E"  ;
    if (arc_index == 147) return "H"  ;
    if (arc_index == 154) return "E"  ;
    if (arc_index == 176) return "W"  ;
    if (arc_index == 178) return "W"  ;
    if (arc_index == 180) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 182) return "W"  ;
    if (arc_index == 184) return "W"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 187) return "W"  ;
    if (arc_index == 188) return "W"  ;
    if (arc_index == 190) return "W"  ;
    if (arc_index == 192) return "W"  ;
    if (arc_index == 193) return "W"  ;
    if (arc_index == 194) return "W"  ;
    if (arc_index == 236) return "H"  ;
    if (arc_index == 250) return "H"  ;
    if (arc_index == 283) return "E"  ;
    if (arc_index == 287) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 304) return "W"  ;
    if (arc_index == 326) return "W"  ;
    if (arc_index == 381) return "H"  ;
    if (arc_index == 413) return "H"  ;
    if (arc_index == 425) return "H"  ;
    if (arc_index == 432) return "H"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 534) return "H"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 620) return "E"  ;
    if (arc_index == 646) return "E"  ;
    if (arc_index == 672) return "E"  ;
    if (arc_index == 685) return "E"  ;
    if (arc_index == 725) return "E"  ;
    if (arc_index == 737) return "E"  ;
    if (arc_index == 741) return "E"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 825) return "W"  ;
    if (arc_index == 871) return "W"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 969) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1035) return "W"  ;
    if (arc_index == 1057) return "E"  ;
    if (arc_index == 1100) return "E"  ;
    if (arc_index == 1124) return "E"  ;
    if (arc_index == 1127) return "W"  ;
    if (arc_index == 1130) return "W"  ;
    if (arc_index == 1136) return "W"  ;
    if (arc_index == 1140) return "W"  ;
    if (arc_index == 1142) return "W"  ;
    if (arc_index == 1173) return "E"  ;
    if (arc_index == 1183) return "H"  ;
    if (arc_index == 1235) return "H"  ;
    if (arc_index == 1239) return "H"  ;
    if (arc_index == 1242) return "H"  ;
    if (arc_index == 1251) return "H"  ;
    if (arc_index == 1253) return "H"  ;
    if (arc_index == 1268) return "H"  ;
    if (arc_index == 1271) return "H"  ;
    if (arc_index == 1278) return "H"  ;
    if (arc_index == 1298) return "H"  ;
    if (arc_index == 1302) return "W"  ;
    if (arc_index == 1304) return "W"  ;
    if (arc_index == 1305) return "W"  ;
    if (arc_index == 1313) return "W"  ;
    if (arc_index == 1316) return "W"  ;
    if (arc_index == 1331) return "W"  ;
    if (arc_index == 1338) return "H"  ;
    if (arc_index == 1342) return "H"  ;
    if (arc_index == 1471) return "H"  ;
    if (arc_index == 1479) return "H"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1566) return "H"  ;
    if (arc_index == 1567) return "H"  ;
    if (arc_index == 1583) return "H"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1686) return "E"  ;
    if (arc_index == 1692) return "H"  ;
    if (arc_index == 1752) return "H"  ;
    if (arc_index == 1770) return "H"  ;
    if (arc_index == 1797) return "E"  ;
    if (arc_index == 1803) return "H"  ;
    if (arc_index == 1836) return "H"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1873) return "H"  ;
    if (arc_index == 1886) return "E"  ;
    if (arc_index == 1900) return "E"  ;
    if (arc_index == 1974) return "E"  ;
    if (arc_index == 2046) return "E"  ;
    if (arc_index == 2048) return "H"  ;
    if (arc_index == 2072) return "H"  ;
    if (arc_index == 2077) return "W"  ;
    if (arc_index == 2079) return "W"  ;
    if (arc_index == 2087) return "W"  ;
    if (arc_index == 2098) return "W"  ;
    if (arc_index == 2130) return "E"  ;
    if (arc_index == 2133) return "E"  ;
    if (arc_index == 2180) return "E"  ;
    if (arc_index == 2195) return "E"  ;
    if (arc_index == 2245) return "H"  ;
    if (arc_index == 2263) return "E"  ;
    if (arc_index == 2288) return "H"  ;
    if (arc_index == 2295) return "H"  ;
    if (arc_index == 2310) return "H"  ;
    if (arc_index == 2311) return "E"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2313) return "W"  ;
    if (arc_index == 2314) return "W"  ;
    if (arc_index == 2315) return "W"  ;
    if (arc_index == 2316) return "W"  ;
    if (arc_index == 2317) return "W"  ;
    if (arc_index == 2318) return "W"  ;
    if (arc_index == 2319) return "W"  ;
    if (arc_index == 2320) return "W"  ;
    if (arc_index == 2321) return "W"  ;
    if (arc_index == 2322) return "W"  ;
    if (arc_index == 2323) return "W"  ;
    if (arc_index == 2324) return "W"  ;
    if (arc_index == 2325) return "W"  ;
    if (arc_index == 2326) return "W"  ;
    if (arc_index == 2327) return "W"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2329) return "W"  ;
    if (arc_index == 2330) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2343) return "H"  ;
    if (arc_index == 2377) return "H"  ;
    if (arc_index == 2388) return "H"  ;
    if (arc_index == 2411) return "W"  ;
    if (arc_index == 2414) return "E"  ;
    if (arc_index == 2444) return "E"  ;
    if (arc_index == 2455) return "E"  ;
    if (arc_index == 2587) return "H"  ;
    if (arc_index == 2594) return "H"  ;
    if (arc_index == 2621) return "H"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2719) return "W"  ;
    if (arc_index == 2725) return "W"  ;
    if (arc_index == 2764) return "H"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2848) return "H"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 9)) begin 
    if (arc_index == 53) return "H"  ;
    if (arc_index == 109) return "E"  ;
    if (arc_index == 124) return "E"  ;
    if (arc_index == 169) return "H"  ;
    if (arc_index == 203) return "H"  ;
    if (arc_index == 243) return "E"  ;
    if (arc_index == 258) return "H"  ;
    if (arc_index == 272) return "H"  ;
    if (arc_index == 300) return "W"  ;
    if (arc_index == 311) return "W"  ;
    if (arc_index == 312) return "W"  ;
    if (arc_index == 315) return "W"  ;
    if (arc_index == 317) return "W"  ;
    if (arc_index == 320) return "W"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 323) return "W"  ;
    if (arc_index == 325) return "W"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 329) return "W"  ;
    if (arc_index == 354) return "E"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 403) return "H"  ;
    if (arc_index == 433) return "H"  ;
    if (arc_index == 536) return "H"  ;
    if (arc_index == 552) return "H"  ;
    if (arc_index == 556) return "H"  ;
    if (arc_index == 558) return "E"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 617) return "W"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 634) return "W"  ;
    if (arc_index == 649) return "E"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 682) return "E"  ;
    if (arc_index == 694) return "E"  ;
    if (arc_index == 713) return "E"  ;
    if (arc_index == 715) return "W"  ;
    if (arc_index == 762) return "E"  ;
    if (arc_index == 820) return "E"  ;
    if (arc_index == 834) return "E"  ;
    if (arc_index == 842) return "E"  ;
    if (arc_index == 846) return "E"  ;
    if (arc_index == 847) return "E"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 1070) return "E"  ;
    if (arc_index == 1142) return "E"  ;
    if (arc_index == 1146) return "E"  ;
    if (arc_index == 1174) return "E"  ;
    if (arc_index == 1205) return "H"  ;
    if (arc_index == 1253) return "H"  ;
    if (arc_index == 1263) return "E"  ;
    if (arc_index == 1323) return "E"  ;
    if (arc_index == 1343) return "E"  ;
    if (arc_index == 1360) return "H"  ;
    if (arc_index == 1379) return "E"  ;
    if (arc_index == 1420) return "E"  ;
    if (arc_index == 1458) return "E"  ;
    if (arc_index == 1493) return "H"  ;
    if (arc_index == 1501) return "H"  ;
    if (arc_index == 1548) return "W"  ;
    if (arc_index == 1558) return "W"  ;
    if (arc_index == 1588) return "H"  ;
    if (arc_index == 1613) return "E"  ;
    if (arc_index == 1714) return "H"  ;
    if (arc_index == 1758) return "H"  ;
    if (arc_index == 1769) return "H"  ;
    if (arc_index == 1770) return "H"  ;
    if (arc_index == 1774) return "H"  ;
    if (arc_index == 1780) return "H"  ;
    if (arc_index == 1825) return "H"  ;
    if (arc_index == 1852) return "H"  ;
    if (arc_index == 1895) return "H"  ;
    if (arc_index == 2068) return "W"  ;
    if (arc_index == 2070) return "H"  ;
    if (arc_index == 2089) return "H"  ;
    if (arc_index == 2092) return "H"  ;
    if (arc_index == 2107) return "E"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2196) return "W"  ;
    if (arc_index == 2262) return "E"  ;
    if (arc_index == 2267) return "H"  ;
    if (arc_index == 2289) return "H"  ;
    if (arc_index == 2310) return "H"  ;
    if (arc_index == 2332) return "H"  ;
    if (arc_index == 2333) return "H"  ;
    if (arc_index == 2334) return "H"  ;
    if (arc_index == 2335) return "W"  ;
    if (arc_index == 2336) return "W"  ;
    if (arc_index == 2337) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2339) return "E"  ;
    if (arc_index == 2340) return "W"  ;
    if (arc_index == 2341) return "W"  ;
    if (arc_index == 2342) return "W"  ;
    if (arc_index == 2343) return "W"  ;
    if (arc_index == 2344) return "W"  ;
    if (arc_index == 2345) return "W"  ;
    if (arc_index == 2346) return "W"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2349) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2351) return "W"  ;
    if (arc_index == 2352) return "W"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2365) return "H"  ;
    if (arc_index == 2380) return "W"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2407) return "W"  ;
    if (arc_index == 2410) return "H"  ;
    if (arc_index == 2467) return "H"  ;
    if (arc_index == 2490) return "E"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2599) return "E"  ;
    if (arc_index == 2600) return "E"  ;
    if (arc_index == 2606) return "E"  ;
    if (arc_index == 2609) return "H"  ;
    if (arc_index == 2611) return "H"  ;
    if (arc_index == 2613) return "H"  ;
    if (arc_index == 2614) return "H"  ;
    if (arc_index == 2615) return "H"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2635) return "W"  ;
    if (arc_index == 2636) return "W"  ;
    if (arc_index == 2637) return "W"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2757) return "E"  ;
    if (arc_index == 2786) return "H"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2870) return "H"  ;
    if (arc_index == 2906) return "W"  ;
    if (arc_index == 2916) return "W"  ;
    if (arc_index == 2923) return "W"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 9)) begin 
    if (arc_index == 17) return "E"  ;
    if (arc_index == 46) return "E"  ;
    if (arc_index == 53) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 75) return "H"  ;
    if (arc_index == 109) return "H"  ;
    if (arc_index == 124) return "H"  ;
    if (arc_index == 168) return "H"  ;
    if (arc_index == 169) return "H"  ;
    if (arc_index == 172) return "E"  ;
    if (arc_index == 191) return "H"  ;
    if (arc_index == 196) return "H"  ;
    if (arc_index == 203) return "E"  ;
    if (arc_index == 213) return "E"  ;
    if (arc_index == 267) return "E"  ;
    if (arc_index == 272) return "E"  ;
    if (arc_index == 280) return "H"  ;
    if (arc_index == 288) return "W"  ;
    if (arc_index == 294) return "H"  ;
    if (arc_index == 301) return "H"  ;
    if (arc_index == 307) return "H"  ;
    if (arc_index == 308) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 321) return "W"  ;
    if (arc_index == 326) return "W"  ;
    if (arc_index == 327) return "W"  ;
    if (arc_index == 400) return "E"  ;
    if (arc_index == 425) return "H"  ;
    if (arc_index == 432) return "H"  ;
    if (arc_index == 526) return "E"  ;
    if (arc_index == 528) return "W"  ;
    if (arc_index == 536) return "W"  ;
    if (arc_index == 566) return "W"  ;
    if (arc_index == 578) return "H"  ;
    if (arc_index == 608) return "W"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 613) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 667) return "W"  ;
    if (arc_index == 685) return "W"  ;
    if (arc_index == 689) return "E"  ;
    if (arc_index == 701) return "E"  ;
    if (arc_index == 706) return "W"  ;
    if (arc_index == 716) return "W"  ;
    if (arc_index == 718) return "W"  ;
    if (arc_index == 792) return "W"  ;
    if (arc_index == 817) return "W"  ;
    if (arc_index == 818) return "W"  ;
    if (arc_index == 823) return "W"  ;
    if (arc_index == 825) return "W"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 829) return "W"  ;
    if (arc_index == 842) return "E"  ;
    if (arc_index == 882) return "E"  ;
    if (arc_index == 975) return "E"  ;
    if (arc_index == 1037) return "E"  ;
    if (arc_index == 1050) return "W"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1103) return "E"  ;
    if (arc_index == 1142) return "E"  ;
    if (arc_index == 1144) return "W"  ;
    if (arc_index == 1145) return "W"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1148) return "W"  ;
    if (arc_index == 1149) return "W"  ;
    if (arc_index == 1150) return "W"  ;
    if (arc_index == 1151) return "W"  ;
    if (arc_index == 1153) return "W"  ;
    if (arc_index == 1156) return "W"  ;
    if (arc_index == 1159) return "W"  ;
    if (arc_index == 1161) return "W"  ;
    if (arc_index == 1162) return "W"  ;
    if (arc_index == 1164) return "W"  ;
    if (arc_index == 1165) return "W"  ;
    if (arc_index == 1177) return "E"  ;
    if (arc_index == 1205) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1227) return "H"  ;
    if (arc_index == 1253) return "H"  ;
    if (arc_index == 1268) return "H"  ;
    if (arc_index == 1316) return "H"  ;
    if (arc_index == 1323) return "H"  ;
    if (arc_index == 1353) return "H"  ;
    if (arc_index == 1356) return "H"  ;
    if (arc_index == 1363) return "H"  ;
    if (arc_index == 1375) return "H"  ;
    if (arc_index == 1382) return "H"  ;
    if (arc_index == 1394) return "H"  ;
    if (arc_index == 1399) return "H"  ;
    if (arc_index == 1421) return "E"  ;
    if (arc_index == 1426) return "E"  ;
    if (arc_index == 1475) return "E"  ;
    if (arc_index == 1515) return "H"  ;
    if (arc_index == 1523) return "H"  ;
    if (arc_index == 1558) return "H"  ;
    if (arc_index == 1577) return "H"  ;
    if (arc_index == 1583) return "H"  ;
    if (arc_index == 1588) return "H"  ;
    if (arc_index == 1598) return "E"  ;
    if (arc_index == 1610) return "H"  ;
    if (arc_index == 1654) return "H"  ;
    if (arc_index == 1680) return "H"  ;
    if (arc_index == 1682) return "E"  ;
    if (arc_index == 1736) return "H"  ;
    if (arc_index == 1769) return "H"  ;
    if (arc_index == 1770) return "H"  ;
    if (arc_index == 1774) return "H"  ;
    if (arc_index == 1780) return "H"  ;
    if (arc_index == 1787) return "E"  ;
    if (arc_index == 1791) return "E"  ;
    if (arc_index == 1797) return "E"  ;
    if (arc_index == 1817) return "E"  ;
    if (arc_index == 1847) return "H"  ;
    if (arc_index == 1869) return "H"  ;
    if (arc_index == 1880) return "H"  ;
    if (arc_index == 1907) return "E"  ;
    if (arc_index == 1917) return "H"  ;
    if (arc_index == 1996) return "E"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2068) return "E"  ;
    if (arc_index == 2070) return "E"  ;
    if (arc_index == 2089) return "E"  ;
    if (arc_index == 2092) return "H"  ;
    if (arc_index == 2100) return "H"  ;
    if (arc_index == 2141) return "E"  ;
    if (arc_index == 2267) return "E"  ;
    if (arc_index == 2286) return "E"  ;
    if (arc_index == 2289) return "H"  ;
    if (arc_index == 2294) return "E"  ;
    if (arc_index == 2295) return "E"  ;
    if (arc_index == 2303) return "E"  ;
    if (arc_index == 2310) return "E"  ;
    if (arc_index == 2326) return "E"  ;
    if (arc_index == 2332) return "H"  ;
    if (arc_index == 2333) return "H"  ;
    if (arc_index == 2336) return "W"  ;
    if (arc_index == 2338) return "W"  ;
    if (arc_index == 2343) return "W"  ;
    if (arc_index == 2345) return "W"  ;
    if (arc_index == 2348) return "W"  ;
    if (arc_index == 2351) return "W"  ;
    if (arc_index == 2354) return "E"  ;
    if (arc_index == 2355) return "W"  ;
    if (arc_index == 2356) return "E"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2358) return "W"  ;
    if (arc_index == 2359) return "W"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2361) return "W"  ;
    if (arc_index == 2362) return "W"  ;
    if (arc_index == 2363) return "W"  ;
    if (arc_index == 2364) return "W"  ;
    if (arc_index == 2365) return "W"  ;
    if (arc_index == 2366) return "W"  ;
    if (arc_index == 2367) return "W"  ;
    if (arc_index == 2368) return "W"  ;
    if (arc_index == 2369) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2371) return "W"  ;
    if (arc_index == 2372) return "W"  ;
    if (arc_index == 2373) return "E"  ;
    if (arc_index == 2374) return "W"  ;
    if (arc_index == 2375) return "W"  ;
    if (arc_index == 2387) return "H"  ;
    if (arc_index == 2403) return "E"  ;
    if (arc_index == 2407) return "E"  ;
    if (arc_index == 2410) return "E"  ;
    if (arc_index == 2415) return "E"  ;
    if (arc_index == 2432) return "H"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2599) return "E"  ;
    if (arc_index == 2606) return "E"  ;
    if (arc_index == 2615) return "E"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2620) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2624) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2627) return "W"  ;
    if (arc_index == 2631) return "H"  ;
    if (arc_index == 2643) return "W"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2775) return "W"  ;
    if (arc_index == 2776) return "W"  ;
    if (arc_index == 2808) return "H"  ;
    if (arc_index == 2830) return "H"  ;
    if (arc_index == 2836) return "H"  ;
    if (arc_index == 2886) return "H"  ;
    if (arc_index == 2892) return "H"  ;
    if (arc_index == 2904) return "H"  ;
    if (arc_index == 2912) return "W"  ;
    if (arc_index == 2922) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 11)) begin 
    if (arc_index == 97) return "H"  ;
    if (arc_index == 146) return "H"  ;
    if (arc_index == 213) return "H"  ;
    if (arc_index == 230) return "H"  ;
    if (arc_index == 302) return "H"  ;
    if (arc_index == 316) return "H"  ;
    if (arc_index == 318) return "H"  ;
    if (arc_index == 447) return "H"  ;
    if (arc_index == 544) return "H"  ;
    if (arc_index == 568) return "H"  ;
    if (arc_index == 600) return "H"  ;
    if (arc_index == 622) return "W"  ;
    if (arc_index == 630) return "W"  ;
    if (arc_index == 632) return "W"  ;
    if (arc_index == 709) return "W"  ;
    if (arc_index == 711) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1050) return "W"  ;
    if (arc_index == 1103) return "W"  ;
    if (arc_index == 1128) return "W"  ;
    if (arc_index == 1249) return "H"  ;
    if (arc_index == 1404) return "H"  ;
    if (arc_index == 1537) return "H"  ;
    if (arc_index == 1545) return "H"  ;
    if (arc_index == 1547) return "H"  ;
    if (arc_index == 1548) return "H"  ;
    if (arc_index == 1552) return "H"  ;
    if (arc_index == 1556) return "H"  ;
    if (arc_index == 1558) return "H"  ;
    if (arc_index == 1632) return "H"  ;
    if (arc_index == 1758) return "H"  ;
    if (arc_index == 1817) return "H"  ;
    if (arc_index == 1869) return "H"  ;
    if (arc_index == 1874) return "H"  ;
    if (arc_index == 1939) return "H"  ;
    if (arc_index == 2073) return "H"  ;
    if (arc_index == 2114) return "H"  ;
    if (arc_index == 2311) return "H"  ;
    if (arc_index == 2354) return "H"  ;
    if (arc_index == 2376) return "W"  ;
    if (arc_index == 2377) return "W"  ;
    if (arc_index == 2378) return "W"  ;
    if (arc_index == 2379) return "W"  ;
    if (arc_index == 2380) return "W"  ;
    if (arc_index == 2381) return "W"  ;
    if (arc_index == 2382) return "W"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2386) return "W"  ;
    if (arc_index == 2387) return "W"  ;
    if (arc_index == 2388) return "W"  ;
    if (arc_index == 2389) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2392) return "W"  ;
    if (arc_index == 2393) return "W"  ;
    if (arc_index == 2394) return "W"  ;
    if (arc_index == 2395) return "W"  ;
    if (arc_index == 2396) return "W"  ;
    if (arc_index == 2397) return "W"  ;
    if (arc_index == 2409) return "H"  ;
    if (arc_index == 2454) return "H"  ;
    if (arc_index == 2618) return "H"  ;
    if (arc_index == 2621) return "H"  ;
    if (arc_index == 2623) return "W"  ;
    if (arc_index == 2632) return "W"  ;
    if (arc_index == 2633) return "W"  ;
    if (arc_index == 2638) return "W"  ;
    if (arc_index == 2639) return "W"  ;
    if (arc_index == 2642) return "W"  ;
    if (arc_index == 2651) return "W"  ;
    if (arc_index == 2653) return "H"  ;
    if (arc_index == 2658) return "H"  ;
    if (arc_index == 2711) return "H"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2727) return "W"  ;
    if (arc_index == 2830) return "H"  ;
    if (arc_index == 2905) return "W"  ;
    if (arc_index == 2907) return "W"  ;
    if (arc_index == 2908) return "W"  ;
    if (arc_index == 2913) return "W"  ;
    if (arc_index == 2914) return "H"  ;
    if (arc_index == 2917) return "H"  ;
    if (arc_index == 2920) return "W"  ;
    if (arc_index == 2921) return "W"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 9)) begin 
    if (arc_index == 8) return "W"  ;
    if (arc_index == 10) return "H"  ;
    if (arc_index == 15) return "E"  ;
    if (arc_index == 24) return "E"  ;
    if (arc_index == 53) return "E"  ;
    if (arc_index == 56) return "E"  ;
    if (arc_index == 75) return "E"  ;
    if (arc_index == 119) return "H"  ;
    if (arc_index == 124) return "H"  ;
    if (arc_index == 168) return "E"  ;
    if (arc_index == 177) return "E"  ;
    if (arc_index == 189) return "E"  ;
    if (arc_index == 193) return "E"  ;
    if (arc_index == 196) return "E"  ;
    if (arc_index == 209) return "E"  ;
    if (arc_index == 221) return "E"  ;
    if (arc_index == 230) return "E"  ;
    if (arc_index == 235) return "H"  ;
    if (arc_index == 250) return "H"  ;
    if (arc_index == 264) return "E"  ;
    if (arc_index == 266) return "E"  ;
    if (arc_index == 293) return "W"  ;
    if (arc_index == 296) return "W"  ;
    if (arc_index == 297) return "W"  ;
    if (arc_index == 299) return "W"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 324) return "H"  ;
    if (arc_index == 326) return "H"  ;
    if (arc_index == 338) return "H"  ;
    if (arc_index == 339) return "H"  ;
    if (arc_index == 341) return "H"  ;
    if (arc_index == 348) return "H"  ;
    if (arc_index == 364) return "E"  ;
    if (arc_index == 413) return "E"  ;
    if (arc_index == 425) return "E"  ;
    if (arc_index == 432) return "E"  ;
    if (arc_index == 447) return "E"  ;
    if (arc_index == 469) return "H"  ;
    if (arc_index == 528) return "H"  ;
    if (arc_index == 529) return "H"  ;
    if (arc_index == 536) return "H"  ;
    if (arc_index == 541) return "W"  ;
    if (arc_index == 545) return "W"  ;
    if (arc_index == 549) return "W"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 596) return "E"  ;
    if (arc_index == 606) return "E"  ;
    if (arc_index == 622) return "H"  ;
    if (arc_index == 636) return "H"  ;
    if (arc_index == 639) return "E"  ;
    if (arc_index == 685) return "E"  ;
    if (arc_index == 704) return "W"  ;
    if (arc_index == 725) return "W"  ;
    if (arc_index == 737) return "W"  ;
    if (arc_index == 741) return "W"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 817) return "E"  ;
    if (arc_index == 818) return "E"  ;
    if (arc_index == 823) return "E"  ;
    if (arc_index == 825) return "E"  ;
    if (arc_index == 922) return "E"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1037) return "E"  ;
    if (arc_index == 1054) return "W"  ;
    if (arc_index == 1066) return "W"  ;
    if (arc_index == 1130) return "W"  ;
    if (arc_index == 1133) return "W"  ;
    if (arc_index == 1136) return "W"  ;
    if (arc_index == 1142) return "W"  ;
    if (arc_index == 1205) return "W"  ;
    if (arc_index == 1242) return "E"  ;
    if (arc_index == 1251) return "E"  ;
    if (arc_index == 1253) return "E"  ;
    if (arc_index == 1255) return "E"  ;
    if (arc_index == 1268) return "E"  ;
    if (arc_index == 1271) return "H"  ;
    if (arc_index == 1277) return "E"  ;
    if (arc_index == 1278) return "E"  ;
    if (arc_index == 1283) return "E"  ;
    if (arc_index == 1298) return "E"  ;
    if (arc_index == 1304) return "W"  ;
    if (arc_index == 1305) return "E"  ;
    if (arc_index == 1313) return "W"  ;
    if (arc_index == 1316) return "W"  ;
    if (arc_index == 1324) return "W"  ;
    if (arc_index == 1331) return "W"  ;
    if (arc_index == 1338) return "W"  ;
    if (arc_index == 1340) return "W"  ;
    if (arc_index == 1361) return "W"  ;
    if (arc_index == 1382) return "W"  ;
    if (arc_index == 1394) return "W"  ;
    if (arc_index == 1399) return "W"  ;
    if (arc_index == 1426) return "H"  ;
    if (arc_index == 1436) return "E"  ;
    if (arc_index == 1479) return "E"  ;
    if (arc_index == 1488) return "E"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1541) return "W"  ;
    if (arc_index == 1542) return "W"  ;
    if (arc_index == 1543) return "W"  ;
    if (arc_index == 1546) return "W"  ;
    if (arc_index == 1549) return "W"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1553) return "W"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1559) return "H"  ;
    if (arc_index == 1567) return "H"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1583) return "W"  ;
    if (arc_index == 1618) return "E"  ;
    if (arc_index == 1654) return "H"  ;
    if (arc_index == 1681) return "E"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1770) return "E"  ;
    if (arc_index == 1780) return "H"  ;
    if (arc_index == 1797) return "H"  ;
    if (arc_index == 1874) return "E"  ;
    if (arc_index == 1880) return "E"  ;
    if (arc_index == 1891) return "H"  ;
    if (arc_index == 1961) return "H"  ;
    if (arc_index == 1975) return "H"  ;
    if (arc_index == 1994) return "E"  ;
    if (arc_index == 2068) return "E"  ;
    if (arc_index == 2070) return "E"  ;
    if (arc_index == 2072) return "W"  ;
    if (arc_index == 2083) return "W"  ;
    if (arc_index == 2100) return "W"  ;
    if (arc_index == 2114) return "E"  ;
    if (arc_index == 2136) return "H"  ;
    if (arc_index == 2141) return "H"  ;
    if (arc_index == 2172) return "H"  ;
    if (arc_index == 2182) return "W"  ;
    if (arc_index == 2186) return "W"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2240) return "E"  ;
    if (arc_index == 2295) return "E"  ;
    if (arc_index == 2310) return "E"  ;
    if (arc_index == 2313) return "W"  ;
    if (arc_index == 2317) return "W"  ;
    if (arc_index == 2320) return "W"  ;
    if (arc_index == 2322) return "W"  ;
    if (arc_index == 2326) return "W"  ;
    if (arc_index == 2329) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2333) return "H"  ;
    if (arc_index == 2343) return "H"  ;
    if (arc_index == 2358) return "E"  ;
    if (arc_index == 2361) return "W"  ;
    if (arc_index == 2376) return "H"  ;
    if (arc_index == 2398) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2400) return "W"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2402) return "W"  ;
    if (arc_index == 2403) return "W"  ;
    if (arc_index == 2404) return "W"  ;
    if (arc_index == 2405) return "W"  ;
    if (arc_index == 2406) return "E"  ;
    if (arc_index == 2407) return "E"  ;
    if (arc_index == 2408) return "E"  ;
    if (arc_index == 2409) return "E"  ;
    if (arc_index == 2410) return "E"  ;
    if (arc_index == 2411) return "E"  ;
    if (arc_index == 2412) return "W"  ;
    if (arc_index == 2413) return "W"  ;
    if (arc_index == 2414) return "W"  ;
    if (arc_index == 2415) return "W"  ;
    if (arc_index == 2416) return "W"  ;
    if (arc_index == 2417) return "W"  ;
    if (arc_index == 2418) return "W"  ;
    if (arc_index == 2419) return "W"  ;
    if (arc_index == 2431) return "H"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2476) return "H"  ;
    if (arc_index == 2482) return "H"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2606) return "E"  ;
    if (arc_index == 2615) return "E"  ;
    if (arc_index == 2623) return "E"  ;
    if (arc_index == 2633) return "E"  ;
    if (arc_index == 2643) return "E"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2675) return "H"  ;
    if (arc_index == 2705) return "E"  ;
    if (arc_index == 2706) return "E"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2714) return "W"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2831) return "E"  ;
    if (arc_index == 2836) return "E"  ;
    if (arc_index == 2852) return "H"  ;
    if (arc_index == 2905) return "H"  ;
    if (arc_index == 2908) return "W"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 3)) begin 
    if (arc_index == 18) return "W"  ;
    if (arc_index == 32) return "H"  ;
    if (arc_index == 42) return "H"  ;
    if (arc_index == 66) return "E"  ;
    if (arc_index == 74) return "E"  ;
    if (arc_index == 141) return "H"  ;
    if (arc_index == 159) return "H"  ;
    if (arc_index == 174) return "H"  ;
    if (arc_index == 186) return "H"  ;
    if (arc_index == 226) return "H"  ;
    if (arc_index == 229) return "H"  ;
    if (arc_index == 238) return "W"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 257) return "H"  ;
    if (arc_index == 268) return "W"  ;
    if (arc_index == 285) return "W"  ;
    if (arc_index == 295) return "W"  ;
    if (arc_index == 346) return "H"  ;
    if (arc_index == 360) return "H"  ;
    if (arc_index == 371) return "W"  ;
    if (arc_index == 386) return "W"  ;
    if (arc_index == 397) return "W"  ;
    if (arc_index == 404) return "W"  ;
    if (arc_index == 405) return "W"  ;
    if (arc_index == 448) return "W"  ;
    if (arc_index == 453) return "E"  ;
    if (arc_index == 461) return "E"  ;
    if (arc_index == 466) return "W"  ;
    if (arc_index == 483) return "W"  ;
    if (arc_index == 488) return "E"  ;
    if (arc_index == 491) return "H"  ;
    if (arc_index == 504) return "E"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 527) return "E"  ;
    if (arc_index == 553) return "E"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 579) return "E"  ;
    if (arc_index == 640) return "W"  ;
    if (arc_index == 644) return "H"  ;
    if (arc_index == 650) return "H"  ;
    if (arc_index == 664) return "H"  ;
    if (arc_index == 668) return "H"  ;
    if (arc_index == 674) return "H"  ;
    if (arc_index == 675) return "H"  ;
    if (arc_index == 676) return "H"  ;
    if (arc_index == 678) return "H"  ;
    if (arc_index == 693) return "H"  ;
    if (arc_index == 703) return "W"  ;
    if (arc_index == 750) return "W"  ;
    if (arc_index == 779) return "E"  ;
    if (arc_index == 802) return "E"  ;
    if (arc_index == 807) return "E"  ;
    if (arc_index == 811) return "E"  ;
    if (arc_index == 858) return "E"  ;
    if (arc_index == 877) return "E"  ;
    if (arc_index == 915) return "E"  ;
    if (arc_index == 928) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 978) return "W"  ;
    if (arc_index == 979) return "W"  ;
    if (arc_index == 993) return "E"  ;
    if (arc_index == 994) return "E"  ;
    if (arc_index == 995) return "E"  ;
    if (arc_index == 996) return "E"  ;
    if (arc_index == 997) return "E"  ;
    if (arc_index == 1000) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1006) return "E"  ;
    if (arc_index == 1008) return "E"  ;
    if (arc_index == 1009) return "E"  ;
    if (arc_index == 1010) return "E"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1027) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1068) return "E"  ;
    if (arc_index == 1131) return "E"  ;
    if (arc_index == 1166) return "W"  ;
    if (arc_index == 1179) return "W"  ;
    if (arc_index == 1184) return "W"  ;
    if (arc_index == 1189) return "E"  ;
    if (arc_index == 1194) return "E"  ;
    if (arc_index == 1195) return "E"  ;
    if (arc_index == 1196) return "E"  ;
    if (arc_index == 1198) return "E"  ;
    if (arc_index == 1199) return "E"  ;
    if (arc_index == 1200) return "E"  ;
    if (arc_index == 1204) return "E"  ;
    if (arc_index == 1206) return "E"  ;
    if (arc_index == 1207) return "E"  ;
    if (arc_index == 1210) return "E"  ;
    if (arc_index == 1211) return "E"  ;
    if (arc_index == 1212) return "E"  ;
    if (arc_index == 1214) return "E"  ;
    if (arc_index == 1215) return "E"  ;
    if (arc_index == 1217) return "E"  ;
    if (arc_index == 1218) return "E"  ;
    if (arc_index == 1222) return "E"  ;
    if (arc_index == 1227) return "E"  ;
    if (arc_index == 1229) return "E"  ;
    if (arc_index == 1230) return "E"  ;
    if (arc_index == 1243) return "W"  ;
    if (arc_index == 1247) return "W"  ;
    if (arc_index == 1266) return "W"  ;
    if (arc_index == 1288) return "W"  ;
    if (arc_index == 1293) return "H"  ;
    if (arc_index == 1318) return "H"  ;
    if (arc_index == 1330) return "W"  ;
    if (arc_index == 1444) return "W"  ;
    if (arc_index == 1448) return "H"  ;
    if (arc_index == 1462) return "W"  ;
    if (arc_index == 1487) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1518) return "E"  ;
    if (arc_index == 1520) return "E"  ;
    if (arc_index == 1521) return "E"  ;
    if (arc_index == 1522) return "E"  ;
    if (arc_index == 1523) return "E"  ;
    if (arc_index == 1525) return "E"  ;
    if (arc_index == 1530) return "E"  ;
    if (arc_index == 1531) return "E"  ;
    if (arc_index == 1537) return "E"  ;
    if (arc_index == 1551) return "W"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1581) return "H"  ;
    if (arc_index == 1589) return "H"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1637) return "E"  ;
    if (arc_index == 1657) return "E"  ;
    if (arc_index == 1658) return "W"  ;
    if (arc_index == 1669) return "W"  ;
    if (arc_index == 1676) return "H"  ;
    if (arc_index == 1723) return "E"  ;
    if (arc_index == 1724) return "E"  ;
    if (arc_index == 1752) return "E"  ;
    if (arc_index == 1753) return "E"  ;
    if (arc_index == 1802) return "H"  ;
    if (arc_index == 1839) return "E"  ;
    if (arc_index == 1842) return "E"  ;
    if (arc_index == 1857) return "W"  ;
    if (arc_index == 1864) return "W"  ;
    if (arc_index == 1913) return "H"  ;
    if (arc_index == 1931) return "H"  ;
    if (arc_index == 1973) return "W"  ;
    if (arc_index == 1983) return "H"  ;
    if (arc_index == 1987) return "H"  ;
    if (arc_index == 2001) return "H"  ;
    if (arc_index == 2006) return "H"  ;
    if (arc_index == 2023) return "H"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2056) return "W"  ;
    if (arc_index == 2062) return "W"  ;
    if (arc_index == 2067) return "W"  ;
    if (arc_index == 2076) return "W"  ;
    if (arc_index == 2134) return "W"  ;
    if (arc_index == 2158) return "H"  ;
    if (arc_index == 2200) return "H"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2227) return "W"  ;
    if (arc_index == 2229) return "E"  ;
    if (arc_index == 2281) return "W"  ;
    if (arc_index == 2312) return "W"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2355) return "H"  ;
    if (arc_index == 2360) return "W"  ;
    if (arc_index == 2370) return "W"  ;
    if (arc_index == 2384) return "W"  ;
    if (arc_index == 2398) return "H"  ;
    if (arc_index == 2420) return "E"  ;
    if (arc_index == 2421) return "E"  ;
    if (arc_index == 2422) return "E"  ;
    if (arc_index == 2423) return "E"  ;
    if (arc_index == 2424) return "E"  ;
    if (arc_index == 2425) return "E"  ;
    if (arc_index == 2426) return "E"  ;
    if (arc_index == 2427) return "E"  ;
    if (arc_index == 2428) return "E"  ;
    if (arc_index == 2429) return "E"  ;
    if (arc_index == 2430) return "E"  ;
    if (arc_index == 2431) return "E"  ;
    if (arc_index == 2432) return "E"  ;
    if (arc_index == 2433) return "E"  ;
    if (arc_index == 2434) return "E"  ;
    if (arc_index == 2435) return "E"  ;
    if (arc_index == 2436) return "W"  ;
    if (arc_index == 2437) return "E"  ;
    if (arc_index == 2438) return "E"  ;
    if (arc_index == 2439) return "E"  ;
    if (arc_index == 2440) return "E"  ;
    if (arc_index == 2441) return "E"  ;
    if (arc_index == 2442) return "E"  ;
    if (arc_index == 2450) return "E"  ;
    if (arc_index == 2452) return "W"  ;
    if (arc_index == 2453) return "H"  ;
    if (arc_index == 2460) return "H"  ;
    if (arc_index == 2483) return "H"  ;
    if (arc_index == 2486) return "H"  ;
    if (arc_index == 2498) return "H"  ;
    if (arc_index == 2508) return "H"  ;
    if (arc_index == 2511) return "E"  ;
    if (arc_index == 2516) return "E"  ;
    if (arc_index == 2540) return "E"  ;
    if (arc_index == 2541) return "E"  ;
    if (arc_index == 2584) return "E"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2672) return "E"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2697) return "H"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2733) return "E"  ;
    if (arc_index == 2755) return "E"  ;
    if (arc_index == 2785) return "E"  ;
    if (arc_index == 2789) return "E"  ;
    if (arc_index == 2796) return "E"  ;
    if (arc_index == 2812) return "E"  ;
    if (arc_index == 2842) return "E"  ;
    if (arc_index == 2854) return "E"  ;
    if (arc_index == 2874) return "H"  ;
    if (arc_index == 2887) return "W"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 4)) begin 
    if (arc_index == 27) return "E"  ;
    if (arc_index == 40) return "E"  ;
    if (arc_index == 48) return "W"  ;
    if (arc_index == 54) return "H"  ;
    if (arc_index == 67) return "H"  ;
    if (arc_index == 110) return "H"  ;
    if (arc_index == 132) return "H"  ;
    if (arc_index == 133) return "H"  ;
    if (arc_index == 135) return "H"  ;
    if (arc_index == 136) return "H"  ;
    if (arc_index == 138) return "H"  ;
    if (arc_index == 142) return "H"  ;
    if (arc_index == 145) return "H"  ;
    if (arc_index == 148) return "H"  ;
    if (arc_index == 149) return "H"  ;
    if (arc_index == 152) return "H"  ;
    if (arc_index == 163) return "H"  ;
    if (arc_index == 165) return "H"  ;
    if (arc_index == 173) return "W"  ;
    if (arc_index == 181) return "W"  ;
    if (arc_index == 210) return "W"  ;
    if (arc_index == 279) return "H"  ;
    if (arc_index == 352) return "H"  ;
    if (arc_index == 355) return "W"  ;
    if (arc_index == 357) return "W"  ;
    if (arc_index == 360) return "W"  ;
    if (arc_index == 368) return "H"  ;
    if (arc_index == 372) return "W"  ;
    if (arc_index == 382) return "H"  ;
    if (arc_index == 392) return "E"  ;
    if (arc_index == 418) return "W"  ;
    if (arc_index == 434) return "W"  ;
    if (arc_index == 439) return "W"  ;
    if (arc_index == 513) return "H"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 638) return "W"  ;
    if (arc_index == 665) return "E"  ;
    if (arc_index == 666) return "H"  ;
    if (arc_index == 669) return "H"  ;
    if (arc_index == 727) return "W"  ;
    if (arc_index == 728) return "W"  ;
    if (arc_index == 732) return "W"  ;
    if (arc_index == 779) return "W"  ;
    if (arc_index == 793) return "E"  ;
    if (arc_index == 795) return "E"  ;
    if (arc_index == 796) return "E"  ;
    if (arc_index == 805) return "E"  ;
    if (arc_index == 806) return "E"  ;
    if (arc_index == 813) return "E"  ;
    if (arc_index == 825) return "W"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 870) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 895) return "W"  ;
    if (arc_index == 927) return "E"  ;
    if (arc_index == 968) return "W"  ;
    if (arc_index == 991) return "E"  ;
    if (arc_index == 992) return "E"  ;
    if (arc_index == 998) return "E"  ;
    if (arc_index == 999) return "E"  ;
    if (arc_index == 1001) return "E"  ;
    if (arc_index == 1003) return "E"  ;
    if (arc_index == 1015) return "E"  ;
    if (arc_index == 1019) return "E"  ;
    if (arc_index == 1031) return "E"  ;
    if (arc_index == 1045) return "E"  ;
    if (arc_index == 1069) return "W"  ;
    if (arc_index == 1123) return "W"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1204) return "E"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1246) return "W"  ;
    if (arc_index == 1267) return "W"  ;
    if (arc_index == 1282) return "W"  ;
    if (arc_index == 1315) return "H"  ;
    if (arc_index == 1371) return "W"  ;
    if (arc_index == 1372) return "W"  ;
    if (arc_index == 1378) return "W"  ;
    if (arc_index == 1381) return "W"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1447) return "W"  ;
    if (arc_index == 1470) return "H"  ;
    if (arc_index == 1496) return "W"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1516) return "W"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1555) return "W"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1603) return "H"  ;
    if (arc_index == 1611) return "H"  ;
    if (arc_index == 1698) return "H"  ;
    if (arc_index == 1724) return "H"  ;
    if (arc_index == 1824) return "H"  ;
    if (arc_index == 1856) return "W"  ;
    if (arc_index == 1931) return "W"  ;
    if (arc_index == 1935) return "H"  ;
    if (arc_index == 1980) return "H"  ;
    if (arc_index == 2005) return "H"  ;
    if (arc_index == 2017) return "E"  ;
    if (arc_index == 2019) return "E"  ;
    if (arc_index == 2137) return "W"  ;
    if (arc_index == 2150) return "E"  ;
    if (arc_index == 2151) return "E"  ;
    if (arc_index == 2164) return "E"  ;
    if (arc_index == 2180) return "H"  ;
    if (arc_index == 2227) return "H"  ;
    if (arc_index == 2279) return "H"  ;
    if (arc_index == 2377) return "H"  ;
    if (arc_index == 2420) return "H"  ;
    if (arc_index == 2442) return "W"  ;
    if (arc_index == 2443) return "W"  ;
    if (arc_index == 2444) return "E"  ;
    if (arc_index == 2445) return "E"  ;
    if (arc_index == 2446) return "E"  ;
    if (arc_index == 2447) return "E"  ;
    if (arc_index == 2448) return "E"  ;
    if (arc_index == 2449) return "E"  ;
    if (arc_index == 2450) return "W"  ;
    if (arc_index == 2451) return "W"  ;
    if (arc_index == 2452) return "W"  ;
    if (arc_index == 2453) return "W"  ;
    if (arc_index == 2454) return "E"  ;
    if (arc_index == 2455) return "E"  ;
    if (arc_index == 2456) return "W"  ;
    if (arc_index == 2457) return "W"  ;
    if (arc_index == 2458) return "W"  ;
    if (arc_index == 2459) return "W"  ;
    if (arc_index == 2460) return "W"  ;
    if (arc_index == 2461) return "W"  ;
    if (arc_index == 2462) return "E"  ;
    if (arc_index == 2463) return "E"  ;
    if (arc_index == 2475) return "H"  ;
    if (arc_index == 2513) return "E"  ;
    if (arc_index == 2514) return "E"  ;
    if (arc_index == 2520) return "H"  ;
    if (arc_index == 2551) return "H"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2577) return "E"  ;
    if (arc_index == 2578) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2592) return "E"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2719) return "H"  ;
    if (arc_index == 2796) return "H"  ;
    if (arc_index == 2812) return "H"  ;
    if (arc_index == 2896) return "H"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 3)) begin 
    if (arc_index == 12) return "W"  ;
    if (arc_index == 26) return "W"  ;
    if (arc_index == 76) return "H"  ;
    if (arc_index == 152) return "W"  ;
    if (arc_index == 185) return "H"  ;
    if (arc_index == 200) return "H"  ;
    if (arc_index == 211) return "W"  ;
    if (arc_index == 244) return "W"  ;
    if (arc_index == 247) return "W"  ;
    if (arc_index == 262) return "W"  ;
    if (arc_index == 301) return "H"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 384) return "E"  ;
    if (arc_index == 390) return "H"  ;
    if (arc_index == 404) return "H"  ;
    if (arc_index == 450) return "H"  ;
    if (arc_index == 472) return "H"  ;
    if (arc_index == 535) return "H"  ;
    if (arc_index == 550) return "W"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 583) return "W"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 664) return "W"  ;
    if (arc_index == 675) return "W"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 688) return "H"  ;
    if (arc_index == 699) return "H"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 751) return "W"  ;
    if (arc_index == 753) return "W"  ;
    if (arc_index == 785) return "W"  ;
    if (arc_index == 815) return "W"  ;
    if (arc_index == 840) return "W"  ;
    if (arc_index == 848) return "W"  ;
    if (arc_index == 849) return "W"  ;
    if (arc_index == 854) return "W"  ;
    if (arc_index == 883) return "E"  ;
    if (arc_index == 887) return "E"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 892) return "E"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 901) return "E"  ;
    if (arc_index == 909) return "E"  ;
    if (arc_index == 914) return "E"  ;
    if (arc_index == 949) return "E"  ;
    if (arc_index == 961) return "E"  ;
    if (arc_index == 1185) return "E"  ;
    if (arc_index == 1193) return "E"  ;
    if (arc_index == 1280) return "E"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1334) return "W"  ;
    if (arc_index == 1337) return "H"  ;
    if (arc_index == 1389) return "H"  ;
    if (arc_index == 1400) return "W"  ;
    if (arc_index == 1407) return "W"  ;
    if (arc_index == 1492) return "H"  ;
    if (arc_index == 1517) return "H"  ;
    if (arc_index == 1587) return "H"  ;
    if (arc_index == 1599) return "E"  ;
    if (arc_index == 1622) return "E"  ;
    if (arc_index == 1625) return "H"  ;
    if (arc_index == 1629) return "H"  ;
    if (arc_index == 1633) return "H"  ;
    if (arc_index == 1667) return "W"  ;
    if (arc_index == 1712) return "W"  ;
    if (arc_index == 1715) return "W"  ;
    if (arc_index == 1718) return "E"  ;
    if (arc_index == 1720) return "H"  ;
    if (arc_index == 1729) return "E"  ;
    if (arc_index == 1739) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1742) return "E"  ;
    if (arc_index == 1747) return "E"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1761) return "E"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1822) return "W"  ;
    if (arc_index == 1828) return "E"  ;
    if (arc_index == 1838) return "E"  ;
    if (arc_index == 1840) return "E"  ;
    if (arc_index == 1846) return "H"  ;
    if (arc_index == 1941) return "H"  ;
    if (arc_index == 1957) return "H"  ;
    if (arc_index == 1959) return "H"  ;
    if (arc_index == 1984) return "W"  ;
    if (arc_index == 1987) return "W"  ;
    if (arc_index == 1993) return "W"  ;
    if (arc_index == 2002) return "W"  ;
    if (arc_index == 2007) return "W"  ;
    if (arc_index == 2024) return "W"  ;
    if (arc_index == 2027) return "H"  ;
    if (arc_index == 2032) return "H"  ;
    if (arc_index == 2034) return "H"  ;
    if (arc_index == 2035) return "H"  ;
    if (arc_index == 2036) return "H"  ;
    if (arc_index == 2038) return "W"  ;
    if (arc_index == 2039) return "W"  ;
    if (arc_index == 2040) return "W"  ;
    if (arc_index == 2042) return "W"  ;
    if (arc_index == 2043) return "W"  ;
    if (arc_index == 2044) return "W"  ;
    if (arc_index == 2050) return "W"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2202) return "H"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2297) return "W"  ;
    if (arc_index == 2399) return "H"  ;
    if (arc_index == 2434) return "E"  ;
    if (arc_index == 2442) return "H"  ;
    if (arc_index == 2464) return "H"  ;
    if (arc_index == 2465) return "E"  ;
    if (arc_index == 2466) return "W"  ;
    if (arc_index == 2467) return "E"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2469) return "E"  ;
    if (arc_index == 2470) return "E"  ;
    if (arc_index == 2471) return "E"  ;
    if (arc_index == 2472) return "E"  ;
    if (arc_index == 2473) return "E"  ;
    if (arc_index == 2474) return "E"  ;
    if (arc_index == 2475) return "E"  ;
    if (arc_index == 2476) return "E"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2478) return "E"  ;
    if (arc_index == 2479) return "W"  ;
    if (arc_index == 2480) return "W"  ;
    if (arc_index == 2481) return "E"  ;
    if (arc_index == 2482) return "E"  ;
    if (arc_index == 2483) return "E"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2485) return "E"  ;
    if (arc_index == 2497) return "H"  ;
    if (arc_index == 2532) return "W"  ;
    if (arc_index == 2542) return "H"  ;
    if (arc_index == 2567) return "H"  ;
    if (arc_index == 2576) return "H"  ;
    if (arc_index == 2597) return "H"  ;
    if (arc_index == 2674) return "H"  ;
    if (arc_index == 2702) return "H"  ;
    if (arc_index == 2706) return "H"  ;
    if (arc_index == 2739) return "H"  ;
    if (arc_index == 2741) return "H"  ;
    if (arc_index == 2743) return "E"  ;
    if (arc_index == 2772) return "W"  ;
    if (arc_index == 2780) return "W"  ;
    if (arc_index == 2788) return "W"  ;
    if (arc_index == 2792) return "W"  ;
    if (arc_index == 2794) return "E"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2801) return "E"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2805) return "E"  ;
    if (arc_index == 2807) return "E"  ;
    if (arc_index == 2810) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2827) return "W"  ;
    if (arc_index == 2840) return "W"  ;
    if (arc_index == 2842) return "W"  ;
    if (arc_index == 2854) return "W"  ;
    if (arc_index == 2856) return "W"  ;
    if (arc_index == 2862) return "E"  ;
    if (arc_index == 2888) return "W"  ;
    if (arc_index == 2893) return "W"  ;
    if (arc_index == 2918) return "H"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 5)) begin 
    if (arc_index == 12) return "H"  ;
    if (arc_index == 14) return "H"  ;
    if (arc_index == 98) return "H"  ;
    if (arc_index == 130) return "H"  ;
    if (arc_index == 142) return "H"  ;
    if (arc_index == 202) return "W"  ;
    if (arc_index == 207) return "H"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 278) return "W"  ;
    if (arc_index == 301) return "W"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 323) return "H"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 367) return "W"  ;
    if (arc_index == 412) return "H"  ;
    if (arc_index == 414) return "H"  ;
    if (arc_index == 426) return "H"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 475) return "E"  ;
    if (arc_index == 480) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 512) return "E"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 553) return "E"  ;
    if (arc_index == 557) return "H"  ;
    if (arc_index == 577) return "H"  ;
    if (arc_index == 611) return "H"  ;
    if (arc_index == 634) return "H"  ;
    if (arc_index == 687) return "H"  ;
    if (arc_index == 690) return "W"  ;
    if (arc_index == 693) return "W"  ;
    if (arc_index == 710) return "H"  ;
    if (arc_index == 717) return "H"  ;
    if (arc_index == 719) return "W"  ;
    if (arc_index == 756) return "E"  ;
    if (arc_index == 757) return "E"  ;
    if (arc_index == 763) return "E"  ;
    if (arc_index == 765) return "E"  ;
    if (arc_index == 784) return "E"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 815) return "E"  ;
    if (arc_index == 816) return "W"  ;
    if (arc_index == 821) return "W"  ;
    if (arc_index == 879) return "W"  ;
    if (arc_index == 883) return "E"  ;
    if (arc_index == 887) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 951) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 967) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1052) return "E"  ;
    if (arc_index == 1062) return "W"  ;
    if (arc_index == 1079) return "W"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1088) return "E"  ;
    if (arc_index == 1089) return "E"  ;
    if (arc_index == 1091) return "E"  ;
    if (arc_index == 1093) return "E"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1149) return "W"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1187) return "W"  ;
    if (arc_index == 1236) return "W"  ;
    if (arc_index == 1257) return "W"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1359) return "H"  ;
    if (arc_index == 1362) return "H"  ;
    if (arc_index == 1390) return "H"  ;
    if (arc_index == 1393) return "H"  ;
    if (arc_index == 1396) return "E"  ;
    if (arc_index == 1397) return "E"  ;
    if (arc_index == 1398) return "E"  ;
    if (arc_index == 1408) return "E"  ;
    if (arc_index == 1411) return "E"  ;
    if (arc_index == 1428) return "E"  ;
    if (arc_index == 1430) return "E"  ;
    if (arc_index == 1432) return "E"  ;
    if (arc_index == 1441) return "E"  ;
    if (arc_index == 1453) return "E"  ;
    if (arc_index == 1455) return "E"  ;
    if (arc_index == 1463) return "E"  ;
    if (arc_index == 1477) return "W"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1484) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1498) return "W"  ;
    if (arc_index == 1514) return "H"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1624) return "E"  ;
    if (arc_index == 1647) return "H"  ;
    if (arc_index == 1655) return "H"  ;
    if (arc_index == 1666) return "E"  ;
    if (arc_index == 1670) return "E"  ;
    if (arc_index == 1672) return "E"  ;
    if (arc_index == 1691) return "E"  ;
    if (arc_index == 1696) return "E"  ;
    if (arc_index == 1698) return "E"  ;
    if (arc_index == 1703) return "E"  ;
    if (arc_index == 1707) return "E"  ;
    if (arc_index == 1710) return "E"  ;
    if (arc_index == 1717) return "E"  ;
    if (arc_index == 1730) return "E"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1736) return "E"  ;
    if (arc_index == 1737) return "E"  ;
    if (arc_index == 1742) return "H"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1751) return "E"  ;
    if (arc_index == 1778) return "W"  ;
    if (arc_index == 1783) return "W"  ;
    if (arc_index == 1784) return "W"  ;
    if (arc_index == 1786) return "W"  ;
    if (arc_index == 1794) return "W"  ;
    if (arc_index == 1798) return "W"  ;
    if (arc_index == 1808) return "W"  ;
    if (arc_index == 1812) return "W"  ;
    if (arc_index == 1826) return "W"  ;
    if (arc_index == 1832) return "E"  ;
    if (arc_index == 1833) return "E"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1837) return "E"  ;
    if (arc_index == 1844) return "E"  ;
    if (arc_index == 1847) return "E"  ;
    if (arc_index == 1852) return "E"  ;
    if (arc_index == 1854) return "E"  ;
    if (arc_index == 1859) return "W"  ;
    if (arc_index == 1862) return "E"  ;
    if (arc_index == 1866) return "E"  ;
    if (arc_index == 1868) return "H"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1895) return "W"  ;
    if (arc_index == 1912) return "W"  ;
    if (arc_index == 1924) return "W"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1958) return "W"  ;
    if (arc_index == 1963) return "W"  ;
    if (arc_index == 1979) return "H"  ;
    if (arc_index == 1982) return "H"  ;
    if (arc_index == 1988) return "H"  ;
    if (arc_index == 1989) return "E"  ;
    if (arc_index == 1991) return "E"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 1996) return "E"  ;
    if (arc_index == 2031) return "E"  ;
    if (arc_index == 2049) return "H"  ;
    if (arc_index == 2055) return "E"  ;
    if (arc_index == 2103) return "W"  ;
    if (arc_index == 2104) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2123) return "E"  ;
    if (arc_index == 2171) return "E"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2224) return "H"  ;
    if (arc_index == 2236) return "E"  ;
    if (arc_index == 2238) return "E"  ;
    if (arc_index == 2257) return "W"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2364) return "W"  ;
    if (arc_index == 2421) return "H"  ;
    if (arc_index == 2464) return "H"  ;
    if (arc_index == 2470) return "E"  ;
    if (arc_index == 2486) return "E"  ;
    if (arc_index == 2487) return "E"  ;
    if (arc_index == 2488) return "W"  ;
    if (arc_index == 2489) return "W"  ;
    if (arc_index == 2490) return "E"  ;
    if (arc_index == 2491) return "E"  ;
    if (arc_index == 2492) return "E"  ;
    if (arc_index == 2493) return "E"  ;
    if (arc_index == 2494) return "E"  ;
    if (arc_index == 2495) return "E"  ;
    if (arc_index == 2496) return "E"  ;
    if (arc_index == 2497) return "W"  ;
    if (arc_index == 2498) return "W"  ;
    if (arc_index == 2499) return "W"  ;
    if (arc_index == 2500) return "W"  ;
    if (arc_index == 2501) return "W"  ;
    if (arc_index == 2502) return "W"  ;
    if (arc_index == 2503) return "E"  ;
    if (arc_index == 2504) return "E"  ;
    if (arc_index == 2505) return "E"  ;
    if (arc_index == 2506) return "E"  ;
    if (arc_index == 2507) return "E"  ;
    if (arc_index == 2519) return "H"  ;
    if (arc_index == 2533) return "H"  ;
    if (arc_index == 2534) return "H"  ;
    if (arc_index == 2535) return "H"  ;
    if (arc_index == 2537) return "H"  ;
    if (arc_index == 2539) return "H"  ;
    if (arc_index == 2540) return "H"  ;
    if (arc_index == 2541) return "H"  ;
    if (arc_index == 2545) return "E"  ;
    if (arc_index == 2549) return "E"  ;
    if (arc_index == 2551) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2564) return "H"  ;
    if (arc_index == 2567) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2603) return "E"  ;
    if (arc_index == 2607) return "E"  ;
    if (arc_index == 2610) return "E"  ;
    if (arc_index == 2627) return "E"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2736) return "W"  ;
    if (arc_index == 2744) return "W"  ;
    if (arc_index == 2749) return "W"  ;
    if (arc_index == 2751) return "E"  ;
    if (arc_index == 2753) return "E"  ;
    if (arc_index == 2763) return "H"  ;
    if (arc_index == 2768) return "E"  ;
    if (arc_index == 2769) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2810) return "E"  ;
    if (arc_index == 2823) return "W"  ;
    if (arc_index == 2827) return "W"  ;
    if (arc_index == 2828) return "W"  ;
    if (arc_index == 2834) return "W"  ;
    if (arc_index == 2835) return "W"  ;
    if (arc_index == 2841) return "W"  ;
    if (arc_index == 2845) return "W"  ;
    if (arc_index == 2849) return "E"  ;
    if (arc_index == 2855) return "E"  ;
    if (arc_index == 2882) return "E"  ;
    if (arc_index == 2901) return "E"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2918) return "W"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 3)) begin 
    if (arc_index == 18) return "W"  ;
    if (arc_index == 36) return "H"  ;
    if (arc_index == 42) return "H"  ;
    if (arc_index == 67) return "E"  ;
    if (arc_index == 93) return "W"  ;
    if (arc_index == 99) return "W"  ;
    if (arc_index == 102) return "W"  ;
    if (arc_index == 112) return "W"  ;
    if (arc_index == 115) return "W"  ;
    if (arc_index == 120) return "H"  ;
    if (arc_index == 135) return "W"  ;
    if (arc_index == 141) return "W"  ;
    if (arc_index == 145) return "W"  ;
    if (arc_index == 159) return "W"  ;
    if (arc_index == 174) return "W"  ;
    if (arc_index == 180) return "W"  ;
    if (arc_index == 186) return "W"  ;
    if (arc_index == 226) return "W"  ;
    if (arc_index == 229) return "H"  ;
    if (arc_index == 246) return "H"  ;
    if (arc_index == 295) return "H"  ;
    if (arc_index == 306) return "W"  ;
    if (arc_index == 345) return "H"  ;
    if (arc_index == 352) return "W"  ;
    if (arc_index == 357) return "W"  ;
    if (arc_index == 360) return "W"  ;
    if (arc_index == 374) return "E"  ;
    if (arc_index == 376) return "E"  ;
    if (arc_index == 377) return "E"  ;
    if (arc_index == 378) return "E"  ;
    if (arc_index == 381) return "E"  ;
    if (arc_index == 382) return "E"  ;
    if (arc_index == 385) return "E"  ;
    if (arc_index == 386) return "E"  ;
    if (arc_index == 387) return "E"  ;
    if (arc_index == 392) return "E"  ;
    if (arc_index == 393) return "E"  ;
    if (arc_index == 397) return "E"  ;
    if (arc_index == 405) return "E"  ;
    if (arc_index == 434) return "H"  ;
    if (arc_index == 448) return "H"  ;
    if (arc_index == 451) return "E"  ;
    if (arc_index == 483) return "E"  ;
    if (arc_index == 524) return "E"  ;
    if (arc_index == 553) return "E"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 579) return "H"  ;
    if (arc_index == 641) return "W"  ;
    if (arc_index == 644) return "W"  ;
    if (arc_index == 645) return "W"  ;
    if (arc_index == 651) return "W"  ;
    if (arc_index == 663) return "E"  ;
    if (arc_index == 664) return "E"  ;
    if (arc_index == 667) return "E"  ;
    if (arc_index == 668) return "E"  ;
    if (arc_index == 674) return "E"  ;
    if (arc_index == 675) return "E"  ;
    if (arc_index == 676) return "E"  ;
    if (arc_index == 678) return "E"  ;
    if (arc_index == 679) return "W"  ;
    if (arc_index == 693) return "W"  ;
    if (arc_index == 732) return "H"  ;
    if (arc_index == 794) return "E"  ;
    if (arc_index == 801) return "E"  ;
    if (arc_index == 807) return "E"  ;
    if (arc_index == 828) return "W"  ;
    if (arc_index == 865) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 915) return "E"  ;
    if (arc_index == 929) return "E"  ;
    if (arc_index == 930) return "E"  ;
    if (arc_index == 933) return "E"  ;
    if (arc_index == 937) return "E"  ;
    if (arc_index == 939) return "E"  ;
    if (arc_index == 940) return "E"  ;
    if (arc_index == 941) return "E"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 993) return "E"  ;
    if (arc_index == 994) return "E"  ;
    if (arc_index == 995) return "E"  ;
    if (arc_index == 996) return "E"  ;
    if (arc_index == 997) return "E"  ;
    if (arc_index == 1000) return "E"  ;
    if (arc_index == 1002) return "W"  ;
    if (arc_index == 1004) return "W"  ;
    if (arc_index == 1005) return "W"  ;
    if (arc_index == 1006) return "W"  ;
    if (arc_index == 1007) return "E"  ;
    if (arc_index == 1008) return "E"  ;
    if (arc_index == 1009) return "E"  ;
    if (arc_index == 1010) return "E"  ;
    if (arc_index == 1014) return "E"  ;
    if (arc_index == 1020) return "E"  ;
    if (arc_index == 1028) return "E"  ;
    if (arc_index == 1033) return "E"  ;
    if (arc_index == 1068) return "E"  ;
    if (arc_index == 1137) return "W"  ;
    if (arc_index == 1198) return "W"  ;
    if (arc_index == 1204) return "E"  ;
    if (arc_index == 1228) return "E"  ;
    if (arc_index == 1240) return "W"  ;
    if (arc_index == 1256) return "W"  ;
    if (arc_index == 1289) return "W"  ;
    if (arc_index == 1371) return "W"  ;
    if (arc_index == 1378) return "W"  ;
    if (arc_index == 1381) return "H"  ;
    if (arc_index == 1439) return "H"  ;
    if (arc_index == 1444) return "H"  ;
    if (arc_index == 1495) return "H"  ;
    if (arc_index == 1496) return "W"  ;
    if (arc_index == 1503) return "W"  ;
    if (arc_index == 1529) return "E"  ;
    if (arc_index == 1536) return "H"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1603) return "E"  ;
    if (arc_index == 1637) return "E"  ;
    if (arc_index == 1657) return "E"  ;
    if (arc_index == 1669) return "H"  ;
    if (arc_index == 1677) return "H"  ;
    if (arc_index == 1687) return "W"  ;
    if (arc_index == 1724) return "E"  ;
    if (arc_index == 1753) return "E"  ;
    if (arc_index == 1764) return "H"  ;
    if (arc_index == 1775) return "H"  ;
    if (arc_index == 1776) return "W"  ;
    if (arc_index == 1842) return "W"  ;
    if (arc_index == 1878) return "W"  ;
    if (arc_index == 1890) return "H"  ;
    if (arc_index == 1931) return "E"  ;
    if (arc_index == 1935) return "E"  ;
    if (arc_index == 1987) return "E"  ;
    if (arc_index == 2001) return "H"  ;
    if (arc_index == 2004) return "E"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2067) return "E"  ;
    if (arc_index == 2071) return "H"  ;
    if (arc_index == 2074) return "W"  ;
    if (arc_index == 2134) return "W"  ;
    if (arc_index == 2140) return "W"  ;
    if (arc_index == 2207) return "W"  ;
    if (arc_index == 2221) return "W"  ;
    if (arc_index == 2227) return "E"  ;
    if (arc_index == 2246) return "H"  ;
    if (arc_index == 2312) return "H"  ;
    if (arc_index == 2328) return "W"  ;
    if (arc_index == 2440) return "W"  ;
    if (arc_index == 2442) return "W"  ;
    if (arc_index == 2443) return "H"  ;
    if (arc_index == 2450) return "H"  ;
    if (arc_index == 2453) return "H"  ;
    if (arc_index == 2461) return "W"  ;
    if (arc_index == 2483) return "E"  ;
    if (arc_index == 2486) return "H"  ;
    if (arc_index == 2508) return "H"  ;
    if (arc_index == 2509) return "H"  ;
    if (arc_index == 2510) return "E"  ;
    if (arc_index == 2511) return "E"  ;
    if (arc_index == 2512) return "E"  ;
    if (arc_index == 2513) return "E"  ;
    if (arc_index == 2514) return "E"  ;
    if (arc_index == 2515) return "W"  ;
    if (arc_index == 2516) return "W"  ;
    if (arc_index == 2517) return "E"  ;
    if (arc_index == 2518) return "E"  ;
    if (arc_index == 2519) return "E"  ;
    if (arc_index == 2520) return "E"  ;
    if (arc_index == 2521) return "E"  ;
    if (arc_index == 2522) return "E"  ;
    if (arc_index == 2523) return "E"  ;
    if (arc_index == 2524) return "E"  ;
    if (arc_index == 2525) return "E"  ;
    if (arc_index == 2526) return "W"  ;
    if (arc_index == 2527) return "W"  ;
    if (arc_index == 2528) return "E"  ;
    if (arc_index == 2529) return "E"  ;
    if (arc_index == 2540) return "E"  ;
    if (arc_index == 2541) return "H"  ;
    if (arc_index == 2586) return "H"  ;
    if (arc_index == 2588) return "E"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2755) return "E"  ;
    if (arc_index == 2785) return "H"  ;
    if (arc_index == 2789) return "H"  ;
    if (arc_index == 2796) return "E"  ;
    if (arc_index == 2842) return "E"  ;
    if (arc_index == 2854) return "W"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 5)) begin 
    if (arc_index == 4) return "W"  ;
    if (arc_index == 12) return "W"  ;
    if (arc_index == 58) return "H"  ;
    if (arc_index == 86) return "H"  ;
    if (arc_index == 130) return "W"  ;
    if (arc_index == 142) return "H"  ;
    if (arc_index == 200) return "W"  ;
    if (arc_index == 204) return "W"  ;
    if (arc_index == 207) return "W"  ;
    if (arc_index == 211) return "W"  ;
    if (arc_index == 244) return "W"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 251) return "H"  ;
    if (arc_index == 273) return "H"  ;
    if (arc_index == 311) return "H"  ;
    if (arc_index == 322) return "W"  ;
    if (arc_index == 323) return "W"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 367) return "H"  ;
    if (arc_index == 414) return "H"  ;
    if (arc_index == 456) return "H"  ;
    if (arc_index == 470) return "H"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 522) return "E"  ;
    if (arc_index == 547) return "E"  ;
    if (arc_index == 550) return "W"  ;
    if (arc_index == 553) return "W"  ;
    if (arc_index == 571) return "W"  ;
    if (arc_index == 574) return "E"  ;
    if (arc_index == 577) return "E"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 601) return "H"  ;
    if (arc_index == 611) return "W"  ;
    if (arc_index == 618) return "W"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 631) return "W"  ;
    if (arc_index == 684) return "W"  ;
    if (arc_index == 687) return "W"  ;
    if (arc_index == 688) return "W"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 699) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 754) return "H"  ;
    if (arc_index == 756) return "H"  ;
    if (arc_index == 757) return "H"  ;
    if (arc_index == 758) return "E"  ;
    if (arc_index == 760) return "E"  ;
    if (arc_index == 762) return "E"  ;
    if (arc_index == 763) return "E"  ;
    if (arc_index == 765) return "E"  ;
    if (arc_index == 771) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 784) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 815) return "W"  ;
    if (arc_index == 826) return "W"  ;
    if (arc_index == 840) return "W"  ;
    if (arc_index == 848) return "W"  ;
    if (arc_index == 849) return "W"  ;
    if (arc_index == 853) return "W"  ;
    if (arc_index == 854) return "W"  ;
    if (arc_index == 879) return "W"  ;
    if (arc_index == 887) return "W"  ;
    if (arc_index == 892) return "E"  ;
    if (arc_index == 893) return "E"  ;
    if (arc_index == 901) return "E"  ;
    if (arc_index == 914) return "E"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 961) return "E"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1076) return "W"  ;
    if (arc_index == 1094) return "E"  ;
    if (arc_index == 1124) return "E"  ;
    if (arc_index == 1187) return "E"  ;
    if (arc_index == 1236) return "W"  ;
    if (arc_index == 1257) return "W"  ;
    if (arc_index == 1321) return "W"  ;
    if (arc_index == 1334) return "W"  ;
    if (arc_index == 1362) return "W"  ;
    if (arc_index == 1390) return "W"  ;
    if (arc_index == 1393) return "W"  ;
    if (arc_index == 1396) return "W"  ;
    if (arc_index == 1397) return "W"  ;
    if (arc_index == 1398) return "W"  ;
    if (arc_index == 1399) return "E"  ;
    if (arc_index == 1401) return "E"  ;
    if (arc_index == 1403) return "H"  ;
    if (arc_index == 1404) return "E"  ;
    if (arc_index == 1405) return "E"  ;
    if (arc_index == 1407) return "W"  ;
    if (arc_index == 1408) return "W"  ;
    if (arc_index == 1411) return "W"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1428) return "W"  ;
    if (arc_index == 1430) return "E"  ;
    if (arc_index == 1432) return "E"  ;
    if (arc_index == 1441) return "E"  ;
    if (arc_index == 1453) return "E"  ;
    if (arc_index == 1463) return "E"  ;
    if (arc_index == 1465) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1473) return "W"  ;
    if (arc_index == 1476) return "W"  ;
    if (arc_index == 1492) return "W"  ;
    if (arc_index == 1498) return "E"  ;
    if (arc_index == 1543) return "W"  ;
    if (arc_index == 1558) return "H"  ;
    if (arc_index == 1599) return "E"  ;
    if (arc_index == 1670) return "E"  ;
    if (arc_index == 1672) return "E"  ;
    if (arc_index == 1691) return "H"  ;
    if (arc_index == 1694) return "W"  ;
    if (arc_index == 1696) return "W"  ;
    if (arc_index == 1697) return "W"  ;
    if (arc_index == 1698) return "W"  ;
    if (arc_index == 1699) return "H"  ;
    if (arc_index == 1702) return "E"  ;
    if (arc_index == 1703) return "E"  ;
    if (arc_index == 1707) return "E"  ;
    if (arc_index == 1710) return "E"  ;
    if (arc_index == 1729) return "E"  ;
    if (arc_index == 1739) return "E"  ;
    if (arc_index == 1742) return "E"  ;
    if (arc_index == 1751) return "E"  ;
    if (arc_index == 1761) return "W"  ;
    if (arc_index == 1768) return "W"  ;
    if (arc_index == 1786) return "H"  ;
    if (arc_index == 1828) return "E"  ;
    if (arc_index == 1833) return "E"  ;
    if (arc_index == 1854) return "E"  ;
    if (arc_index == 1866) return "E"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1895) return "E"  ;
    if (arc_index == 1912) return "H"  ;
    if (arc_index == 1924) return "H"  ;
    if (arc_index == 1959) return "W"  ;
    if (arc_index == 1985) return "E"  ;
    if (arc_index == 1986) return "E"  ;
    if (arc_index == 1988) return "E"  ;
    if (arc_index == 1989) return "E"  ;
    if (arc_index == 1990) return "E"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 1997) return "E"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2023) return "H"  ;
    if (arc_index == 2031) return "H"  ;
    if (arc_index == 2093) return "H"  ;
    if (arc_index == 2096) return "W"  ;
    if (arc_index == 2104) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2192) return "W"  ;
    if (arc_index == 2223) return "W"  ;
    if (arc_index == 2238) return "W"  ;
    if (arc_index == 2265) return "W"  ;
    if (arc_index == 2268) return "H"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2465) return "H"  ;
    if (arc_index == 2467) return "E"  ;
    if (arc_index == 2468) return "E"  ;
    if (arc_index == 2471) return "E"  ;
    if (arc_index == 2476) return "E"  ;
    if (arc_index == 2481) return "E"  ;
    if (arc_index == 2482) return "E"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2487) return "E"  ;
    if (arc_index == 2501) return "E"  ;
    if (arc_index == 2508) return "H"  ;
    if (arc_index == 2530) return "H"  ;
    if (arc_index == 2531) return "E"  ;
    if (arc_index == 2532) return "W"  ;
    if (arc_index == 2533) return "W"  ;
    if (arc_index == 2534) return "W"  ;
    if (arc_index == 2535) return "W"  ;
    if (arc_index == 2536) return "W"  ;
    if (arc_index == 2537) return "W"  ;
    if (arc_index == 2538) return "E"  ;
    if (arc_index == 2539) return "E"  ;
    if (arc_index == 2540) return "E"  ;
    if (arc_index == 2541) return "E"  ;
    if (arc_index == 2542) return "W"  ;
    if (arc_index == 2543) return "E"  ;
    if (arc_index == 2544) return "E"  ;
    if (arc_index == 2545) return "E"  ;
    if (arc_index == 2546) return "E"  ;
    if (arc_index == 2547) return "W"  ;
    if (arc_index == 2548) return "E"  ;
    if (arc_index == 2549) return "E"  ;
    if (arc_index == 2550) return "E"  ;
    if (arc_index == 2551) return "E"  ;
    if (arc_index == 2554) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2563) return "H"  ;
    if (arc_index == 2564) return "H"  ;
    if (arc_index == 2573) return "H"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2603) return "E"  ;
    if (arc_index == 2607) return "E"  ;
    if (arc_index == 2608) return "H"  ;
    if (arc_index == 2627) return "W"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2736) return "W"  ;
    if (arc_index == 2744) return "W"  ;
    if (arc_index == 2749) return "W"  ;
    if (arc_index == 2757) return "E"  ;
    if (arc_index == 2779) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2786) return "E"  ;
    if (arc_index == 2790) return "E"  ;
    if (arc_index == 2794) return "E"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2807) return "H"  ;
    if (arc_index == 2810) return "H"  ;
    if (arc_index == 2832) return "W"  ;
    if (arc_index == 2835) return "W"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2841) return "E"  ;
    if (arc_index == 2845) return "E"  ;
    if (arc_index == 2849) return "E"  ;
    if (arc_index == 2862) return "E"  ;
    if (arc_index == 2918) return "W"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 1)) begin 
    if (arc_index == 80) return "H"  ;
    if (arc_index == 164) return "H"  ;
    if (arc_index == 273) return "H"  ;
    if (arc_index == 389) return "H"  ;
    if (arc_index == 478) return "H"  ;
    if (arc_index == 492) return "H"  ;
    if (arc_index == 565) return "H"  ;
    if (arc_index == 623) return "H"  ;
    if (arc_index == 773) return "H"  ;
    if (arc_index == 776) return "H"  ;
    if (arc_index == 786) return "W"  ;
    if (arc_index == 1425) return "H"  ;
    if (arc_index == 1580) return "H"  ;
    if (arc_index == 1713) return "H"  ;
    if (arc_index == 1721) return "H"  ;
    if (arc_index == 1808) return "H"  ;
    if (arc_index == 1934) return "H"  ;
    if (arc_index == 2045) return "H"  ;
    if (arc_index == 2110) return "H"  ;
    if (arc_index == 2115) return "H"  ;
    if (arc_index == 2290) return "H"  ;
    if (arc_index == 2487) return "H"  ;
    if (arc_index == 2530) return "H"  ;
    if (arc_index == 2552) return "H"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2554) return "E"  ;
    if (arc_index == 2555) return "E"  ;
    if (arc_index == 2556) return "E"  ;
    if (arc_index == 2557) return "E"  ;
    if (arc_index == 2558) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2560) return "E"  ;
    if (arc_index == 2561) return "E"  ;
    if (arc_index == 2562) return "E"  ;
    if (arc_index == 2563) return "E"  ;
    if (arc_index == 2564) return "E"  ;
    if (arc_index == 2565) return "E"  ;
    if (arc_index == 2566) return "E"  ;
    if (arc_index == 2567) return "E"  ;
    if (arc_index == 2568) return "E"  ;
    if (arc_index == 2569) return "E"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2571) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2585) return "H"  ;
    if (arc_index == 2630) return "H"  ;
    if (arc_index == 2829) return "H"  ;
    if (arc_index == 2859) return "H"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 1)) begin 
    if (arc_index == 102) return "H"  ;
    if (arc_index == 186) return "H"  ;
    if (arc_index == 268) return "H"  ;
    if (arc_index == 295) return "H"  ;
    if (arc_index == 394) return "H"  ;
    if (arc_index == 407) return "H"  ;
    if (arc_index == 411) return "H"  ;
    if (arc_index == 418) return "H"  ;
    if (arc_index == 500) return "H"  ;
    if (arc_index == 505) return "H"  ;
    if (arc_index == 514) return "H"  ;
    if (arc_index == 575) return "H"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 645) return "H"  ;
    if (arc_index == 750) return "H"  ;
    if (arc_index == 798) return "H"  ;
    if (arc_index == 947) return "H"  ;
    if (arc_index == 1013) return "H"  ;
    if (arc_index == 1016) return "H"  ;
    if (arc_index == 1017) return "H"  ;
    if (arc_index == 1018) return "H"  ;
    if (arc_index == 1020) return "H"  ;
    if (arc_index == 1021) return "H"  ;
    if (arc_index == 1022) return "H"  ;
    if (arc_index == 1024) return "H"  ;
    if (arc_index == 1025) return "H"  ;
    if (arc_index == 1026) return "H"  ;
    if (arc_index == 1027) return "H"  ;
    if (arc_index == 1028) return "H"  ;
    if (arc_index == 1029) return "H"  ;
    if (arc_index == 1032) return "H"  ;
    if (arc_index == 1090) return "H"  ;
    if (arc_index == 1447) return "H"  ;
    if (arc_index == 1466) return "H"  ;
    if (arc_index == 1526) return "H"  ;
    if (arc_index == 1602) return "H"  ;
    if (arc_index == 1659) return "H"  ;
    if (arc_index == 1735) return "H"  ;
    if (arc_index == 1743) return "H"  ;
    if (arc_index == 1830) return "H"  ;
    if (arc_index == 1864) return "H"  ;
    if (arc_index == 1878) return "H"  ;
    if (arc_index == 1956) return "H"  ;
    if (arc_index == 2067) return "H"  ;
    if (arc_index == 2137) return "H"  ;
    if (arc_index == 2162) return "H"  ;
    if (arc_index == 2230) return "E"  ;
    if (arc_index == 2312) return "H"  ;
    if (arc_index == 2509) return "H"  ;
    if (arc_index == 2552) return "H"  ;
    if (arc_index == 2574) return "H"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2576) return "E"  ;
    if (arc_index == 2577) return "E"  ;
    if (arc_index == 2578) return "E"  ;
    if (arc_index == 2579) return "E"  ;
    if (arc_index == 2580) return "E"  ;
    if (arc_index == 2581) return "E"  ;
    if (arc_index == 2582) return "E"  ;
    if (arc_index == 2583) return "E"  ;
    if (arc_index == 2584) return "E"  ;
    if (arc_index == 2585) return "E"  ;
    if (arc_index == 2586) return "E"  ;
    if (arc_index == 2587) return "E"  ;
    if (arc_index == 2588) return "E"  ;
    if (arc_index == 2589) return "E"  ;
    if (arc_index == 2590) return "E"  ;
    if (arc_index == 2591) return "E"  ;
    if (arc_index == 2592) return "E"  ;
    if (arc_index == 2593) return "E"  ;
    if (arc_index == 2594) return "E"  ;
    if (arc_index == 2595) return "E"  ;
    if (arc_index == 2607) return "H"  ;
    if (arc_index == 2652) return "H"  ;
    if (arc_index == 2811) return "H"  ;
    if (arc_index == 2851) return "H"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 9)) begin 
    if (arc_index == 86) return "E"  ;
    if (arc_index == 124) return "H"  ;
    if (arc_index == 208) return "H"  ;
    if (arc_index == 243) return "H"  ;
    if (arc_index == 254) return "E"  ;
    if (arc_index == 258) return "E"  ;
    if (arc_index == 317) return "H"  ;
    if (arc_index == 433) return "H"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 522) return "H"  ;
    if (arc_index == 536) return "H"  ;
    if (arc_index == 558) return "H"  ;
    if (arc_index == 563) return "E"  ;
    if (arc_index == 621) return "W"  ;
    if (arc_index == 667) return "H"  ;
    if (arc_index == 682) return "E"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 708) return "W"  ;
    if (arc_index == 710) return "W"  ;
    if (arc_index == 712) return "W"  ;
    if (arc_index == 713) return "W"  ;
    if (arc_index == 715) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 719) return "W"  ;
    if (arc_index == 720) return "W"  ;
    if (arc_index == 721) return "W"  ;
    if (arc_index == 722) return "W"  ;
    if (arc_index == 782) return "E"  ;
    if (arc_index == 820) return "H"  ;
    if (arc_index == 834) return "W"  ;
    if (arc_index == 1142) return "W"  ;
    if (arc_index == 1146) return "W"  ;
    if (arc_index == 1253) return "W"  ;
    if (arc_index == 1323) return "W"  ;
    if (arc_index == 1343) return "W"  ;
    if (arc_index == 1467) return "E"  ;
    if (arc_index == 1468) return "E"  ;
    if (arc_index == 1469) return "H"  ;
    if (arc_index == 1547) return "H"  ;
    if (arc_index == 1624) return "H"  ;
    if (arc_index == 1701) return "E"  ;
    if (arc_index == 1757) return "H"  ;
    if (arc_index == 1758) return "H"  ;
    if (arc_index == 1765) return "H"  ;
    if (arc_index == 1769) return "H"  ;
    if (arc_index == 1770) return "H"  ;
    if (arc_index == 1774) return "H"  ;
    if (arc_index == 1780) return "H"  ;
    if (arc_index == 1852) return "H"  ;
    if (arc_index == 1854) return "E"  ;
    if (arc_index == 1978) return "H"  ;
    if (arc_index == 2089) return "H"  ;
    if (arc_index == 2092) return "H"  ;
    if (arc_index == 2107) return "H"  ;
    if (arc_index == 2159) return "H"  ;
    if (arc_index == 2289) return "H"  ;
    if (arc_index == 2334) return "H"  ;
    if (arc_index == 2337) return "W"  ;
    if (arc_index == 2349) return "W"  ;
    if (arc_index == 2407) return "W"  ;
    if (arc_index == 2503) return "E"  ;
    if (arc_index == 2531) return "H"  ;
    if (arc_index == 2574) return "H"  ;
    if (arc_index == 2596) return "E"  ;
    if (arc_index == 2597) return "W"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2599) return "W"  ;
    if (arc_index == 2600) return "W"  ;
    if (arc_index == 2601) return "W"  ;
    if (arc_index == 2602) return "W"  ;
    if (arc_index == 2603) return "W"  ;
    if (arc_index == 2604) return "W"  ;
    if (arc_index == 2605) return "W"  ;
    if (arc_index == 2606) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2608) return "W"  ;
    if (arc_index == 2609) return "W"  ;
    if (arc_index == 2610) return "W"  ;
    if (arc_index == 2611) return "W"  ;
    if (arc_index == 2612) return "W"  ;
    if (arc_index == 2613) return "W"  ;
    if (arc_index == 2614) return "W"  ;
    if (arc_index == 2615) return "W"  ;
    if (arc_index == 2616) return "E"  ;
    if (arc_index == 2617) return "W"  ;
    if (arc_index == 2626) return "W"  ;
    if (arc_index == 2629) return "H"  ;
    if (arc_index == 2674) return "H"  ;
    if (arc_index == 2757) return "H"  ;
    if (arc_index == 2791) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2873) return "H"  ;
  end 
  if ((thisRowAddr == 4) & (thisColAddr == 11)) begin 
    if (arc_index == 146) return "H"  ;
    if (arc_index == 179) return "H"  ;
    if (arc_index == 230) return "H"  ;
    if (arc_index == 318) return "H"  ;
    if (arc_index == 339) return "H"  ;
    if (arc_index == 455) return "H"  ;
    if (arc_index == 544) return "H"  ;
    if (arc_index == 558) return "H"  ;
    if (arc_index == 568) return "H"  ;
    if (arc_index == 616) return "W"  ;
    if (arc_index == 620) return "W"  ;
    if (arc_index == 622) return "W"  ;
    if (arc_index == 626) return "W"  ;
    if (arc_index == 630) return "W"  ;
    if (arc_index == 632) return "W"  ;
    if (arc_index == 636) return "W"  ;
    if (arc_index == 637) return "W"  ;
    if (arc_index == 689) return "H"  ;
    if (arc_index == 709) return "H"  ;
    if (arc_index == 711) return "H"  ;
    if (arc_index == 741) return "H"  ;
    if (arc_index == 842) return "H"  ;
    if (arc_index == 1103) return "H"  ;
    if (arc_index == 1128) return "H"  ;
    if (arc_index == 1404) return "H"  ;
    if (arc_index == 1491) return "H"  ;
    if (arc_index == 1547) return "H"  ;
    if (arc_index == 1548) return "H"  ;
    if (arc_index == 1552) return "W"  ;
    if (arc_index == 1556) return "W"  ;
    if (arc_index == 1558) return "W"  ;
    if (arc_index == 1646) return "H"  ;
    if (arc_index == 1758) return "H"  ;
    if (arc_index == 1779) return "H"  ;
    if (arc_index == 1787) return "H"  ;
    if (arc_index == 1817) return "H"  ;
    if (arc_index == 1874) return "H"  ;
    if (arc_index == 2000) return "H"  ;
    if (arc_index == 2073) return "H"  ;
    if (arc_index == 2111) return "H"  ;
    if (arc_index == 2181) return "H"  ;
    if (arc_index == 2356) return "H"  ;
    if (arc_index == 2379) return "H"  ;
    if (arc_index == 2380) return "H"  ;
    if (arc_index == 2383) return "H"  ;
    if (arc_index == 2385) return "H"  ;
    if (arc_index == 2397) return "H"  ;
    if (arc_index == 2415) return "H"  ;
    if (arc_index == 2553) return "H"  ;
    if (arc_index == 2596) return "H"  ;
    if (arc_index == 2618) return "H"  ;
    if (arc_index == 2619) return "W"  ;
    if (arc_index == 2620) return "W"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2622) return "W"  ;
    if (arc_index == 2623) return "W"  ;
    if (arc_index == 2624) return "W"  ;
    if (arc_index == 2625) return "W"  ;
    if (arc_index == 2626) return "W"  ;
    if (arc_index == 2627) return "W"  ;
    if (arc_index == 2628) return "W"  ;
    if (arc_index == 2629) return "W"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2631) return "W"  ;
    if (arc_index == 2632) return "W"  ;
    if (arc_index == 2633) return "W"  ;
    if (arc_index == 2634) return "W"  ;
    if (arc_index == 2635) return "W"  ;
    if (arc_index == 2636) return "W"  ;
    if (arc_index == 2637) return "W"  ;
    if (arc_index == 2638) return "W"  ;
    if (arc_index == 2639) return "W"  ;
    if (arc_index == 2642) return "W"  ;
    if (arc_index == 2651) return "H"  ;
    if (arc_index == 2658) return "H"  ;
    if (arc_index == 2696) return "H"  ;
    if (arc_index == 2711) return "H"  ;
    if (arc_index == 2895) return "H"  ;
    if (arc_index == 2905) return "H"  ;
    if (arc_index == 2907) return "H"  ;
    if (arc_index == 2908) return "H"  ;
    if (arc_index == 2913) return "H"  ;
    if (arc_index == 2914) return "H"  ;
    if (arc_index == 2917) return "H"  ;
    if (arc_index == 2920) return "H"  ;
    if (arc_index == 2921) return "H"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 11)) begin 
    if (arc_index == 168) return "H"  ;
    if (arc_index == 252) return "H"  ;
    if (arc_index == 361) return "H"  ;
    if (arc_index == 477) return "H"  ;
    if (arc_index == 566) return "H"  ;
    if (arc_index == 580) return "H"  ;
    if (arc_index == 711) return "H"  ;
    if (arc_index == 864) return "H"  ;
    if (arc_index == 1513) return "H"  ;
    if (arc_index == 1668) return "H"  ;
    if (arc_index == 1801) return "H"  ;
    if (arc_index == 1809) return "H"  ;
    if (arc_index == 1896) return "H"  ;
    if (arc_index == 2022) return "H"  ;
    if (arc_index == 2133) return "H"  ;
    if (arc_index == 2203) return "H"  ;
    if (arc_index == 2378) return "H"  ;
    if (arc_index == 2575) return "H"  ;
    if (arc_index == 2618) return "H"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2641) return "W"  ;
    if (arc_index == 2642) return "W"  ;
    if (arc_index == 2643) return "W"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2646) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2650) return "W"  ;
    if (arc_index == 2651) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2653) return "W"  ;
    if (arc_index == 2654) return "W"  ;
    if (arc_index == 2655) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2657) return "W"  ;
    if (arc_index == 2658) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2660) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2673) return "H"  ;
    if (arc_index == 2718) return "H"  ;
    if (arc_index == 2917) return "H"  ;
  end 
  if ((thisRowAddr == 6) & (thisColAddr == 0)) begin 
    if (arc_index == 13) return "H"  ;
    if (arc_index == 135) return "H"  ;
    if (arc_index == 190) return "H"  ;
    if (arc_index == 274) return "H"  ;
    if (arc_index == 383) return "H"  ;
    if (arc_index == 388) return "H"  ;
    if (arc_index == 457) return "H"  ;
    if (arc_index == 485) return "H"  ;
    if (arc_index == 486) return "H"  ;
    if (arc_index == 492) return "H"  ;
    if (arc_index == 493) return "H"  ;
    if (arc_index == 494) return "H"  ;
    if (arc_index == 499) return "H"  ;
    if (arc_index == 503) return "H"  ;
    if (arc_index == 573) return "E"  ;
    if (arc_index == 575) return "E"  ;
    if (arc_index == 579) return "E"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 582) return "E"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 588) return "H"  ;
    if (arc_index == 592) return "H"  ;
    if (arc_index == 602) return "H"  ;
    if (arc_index == 733) return "H"  ;
    if (arc_index == 761) return "H"  ;
    if (arc_index == 774) return "H"  ;
    if (arc_index == 886) return "H"  ;
    if (arc_index == 947) return "H"  ;
    if (arc_index == 957) return "E"  ;
    if (arc_index == 1026) return "E"  ;
    if (arc_index == 1081) return "E"  ;
    if (arc_index == 1219) return "E"  ;
    if (arc_index == 1453) return "E"  ;
    if (arc_index == 1481) return "E"  ;
    if (arc_index == 1519) return "E"  ;
    if (arc_index == 1532) return "E"  ;
    if (arc_index == 1534) return "E"  ;
    if (arc_index == 1535) return "H"  ;
    if (arc_index == 1562) return "H"  ;
    if (arc_index == 1589) return "H"  ;
    if (arc_index == 1590) return "E"  ;
    if (arc_index == 1592) return "E"  ;
    if (arc_index == 1596) return "E"  ;
    if (arc_index == 1602) return "E"  ;
    if (arc_index == 1603) return "E"  ;
    if (arc_index == 1690) return "H"  ;
    if (arc_index == 1823) return "H"  ;
    if (arc_index == 1831) return "H"  ;
    if (arc_index == 1918) return "H"  ;
    if (arc_index == 2044) return "H"  ;
    if (arc_index == 2155) return "H"  ;
    if (arc_index == 2225) return "H"  ;
    if (arc_index == 2231) return "H"  ;
    if (arc_index == 2400) return "H"  ;
    if (arc_index == 2436) return "H"  ;
    if (arc_index == 2571) return "H"  ;
    if (arc_index == 2581) return "H"  ;
    if (arc_index == 2597) return "H"  ;
    if (arc_index == 2640) return "H"  ;
    if (arc_index == 2662) return "E"  ;
    if (arc_index == 2663) return "E"  ;
    if (arc_index == 2664) return "E"  ;
    if (arc_index == 2665) return "E"  ;
    if (arc_index == 2666) return "E"  ;
    if (arc_index == 2667) return "E"  ;
    if (arc_index == 2668) return "E"  ;
    if (arc_index == 2669) return "E"  ;
    if (arc_index == 2670) return "E"  ;
    if (arc_index == 2671) return "E"  ;
    if (arc_index == 2672) return "E"  ;
    if (arc_index == 2673) return "E"  ;
    if (arc_index == 2674) return "E"  ;
    if (arc_index == 2675) return "E"  ;
    if (arc_index == 2676) return "E"  ;
    if (arc_index == 2677) return "E"  ;
    if (arc_index == 2678) return "E"  ;
    if (arc_index == 2679) return "E"  ;
    if (arc_index == 2680) return "E"  ;
    if (arc_index == 2681) return "E"  ;
    if (arc_index == 2682) return "E"  ;
    if (arc_index == 2683) return "E"  ;
    if (arc_index == 2695) return "H"  ;
    if (arc_index == 2740) return "H"  ;
    if (arc_index == 2792) return "H"  ;
    if (arc_index == 2874) return "E"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2879) return "E"  ;
    if (arc_index == 2903) return "E"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 3)) begin 
    if (arc_index == 7) return "W"  ;
    if (arc_index == 13) return "W"  ;
    if (arc_index == 18) return "W"  ;
    if (arc_index == 35) return "H"  ;
    if (arc_index == 41) return "H"  ;
    if (arc_index == 49) return "H"  ;
    if (arc_index == 50) return "H"  ;
    if (arc_index == 76) return "H"  ;
    if (arc_index == 152) return "H"  ;
    if (arc_index == 158) return "H"  ;
    if (arc_index == 160) return "W"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 200) return "W"  ;
    if (arc_index == 212) return "H"  ;
    if (arc_index == 246) return "H"  ;
    if (arc_index == 296) return "H"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 404) return "W"  ;
    if (arc_index == 405) return "H"  ;
    if (arc_index == 406) return "W"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 454) return "E"  ;
    if (arc_index == 470) return "E"  ;
    if (arc_index == 471) return "E"  ;
    if (arc_index == 472) return "E"  ;
    if (arc_index == 475) return "E"  ;
    if (arc_index == 478) return "E"  ;
    if (arc_index == 479) return "E"  ;
    if (arc_index == 480) return "E"  ;
    if (arc_index == 482) return "E"  ;
    if (arc_index == 494) return "E"  ;
    if (arc_index == 506) return "E"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 521) return "H"  ;
    if (arc_index == 524) return "H"  ;
    if (arc_index == 525) return "H"  ;
    if (arc_index == 553) return "H"  ;
    if (arc_index == 570) return "H"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 602) return "E"  ;
    if (arc_index == 610) return "H"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 624) return "H"  ;
    if (arc_index == 650) return "W"  ;
    if (arc_index == 654) return "W"  ;
    if (arc_index == 656) return "W"  ;
    if (arc_index == 664) return "W"  ;
    if (arc_index == 675) return "W"  ;
    if (arc_index == 676) return "E"  ;
    if (arc_index == 678) return "E"  ;
    if (arc_index == 693) return "E"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 734) return "W"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 750) return "W"  ;
    if (arc_index == 755) return "H"  ;
    if (arc_index == 785) return "E"  ;
    if (arc_index == 808) return "E"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 811) return "E"  ;
    if (arc_index == 858) return "W"  ;
    if (arc_index == 877) return "W"  ;
    if (arc_index == 888) return "W"  ;
    if (arc_index == 890) return "E"  ;
    if (arc_index == 895) return "E"  ;
    if (arc_index == 896) return "E"  ;
    if (arc_index == 898) return "E"  ;
    if (arc_index == 908) return "H"  ;
    if (arc_index == 914) return "H"  ;
    if (arc_index == 921) return "H"  ;
    if (arc_index == 953) return "E"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 956) return "E"  ;
    if (arc_index == 987) return "E"  ;
    if (arc_index == 994) return "E"  ;
    if (arc_index == 995) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1032) return "E"  ;
    if (arc_index == 1044) return "E"  ;
    if (arc_index == 1063) return "E"  ;
    if (arc_index == 1075) return "W"  ;
    if (arc_index == 1077) return "W"  ;
    if (arc_index == 1096) return "W"  ;
    if (arc_index == 1121) return "W"  ;
    if (arc_index == 1143) return "W"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1170) return "W"  ;
    if (arc_index == 1190) return "E"  ;
    if (arc_index == 1208) return "E"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1269) return "E"  ;
    if (arc_index == 1279) return "E"  ;
    if (arc_index == 1296) return "W"  ;
    if (arc_index == 1301) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1459) return "W"  ;
    if (arc_index == 1465) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1557) return "H"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1594) return "E"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1599) return "E"  ;
    if (arc_index == 1606) return "W"  ;
    if (arc_index == 1612) return "W"  ;
    if (arc_index == 1617) return "W"  ;
    if (arc_index == 1629) return "W"  ;
    if (arc_index == 1630) return "E"  ;
    if (arc_index == 1631) return "E"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1633) return "E"  ;
    if (arc_index == 1635) return "E"  ;
    if (arc_index == 1638) return "E"  ;
    if (arc_index == 1639) return "E"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1641) return "E"  ;
    if (arc_index == 1645) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1648) return "E"  ;
    if (arc_index == 1649) return "E"  ;
    if (arc_index == 1657) return "E"  ;
    if (arc_index == 1658) return "E"  ;
    if (arc_index == 1659) return "E"  ;
    if (arc_index == 1660) return "E"  ;
    if (arc_index == 1669) return "E"  ;
    if (arc_index == 1674) return "W"  ;
    if (arc_index == 1683) return "W"  ;
    if (arc_index == 1712) return "H"  ;
    if (arc_index == 1715) return "H"  ;
    if (arc_index == 1724) return "H"  ;
    if (arc_index == 1731) return "E"  ;
    if (arc_index == 1753) return "E"  ;
    if (arc_index == 1790) return "E"  ;
    if (arc_index == 1795) return "E"  ;
    if (arc_index == 1823) return "E"  ;
    if (arc_index == 1827) return "E"  ;
    if (arc_index == 1834) return "E"  ;
    if (arc_index == 1835) return "W"  ;
    if (arc_index == 1839) return "W"  ;
    if (arc_index == 1842) return "W"  ;
    if (arc_index == 1843) return "W"  ;
    if (arc_index == 1845) return "H"  ;
    if (arc_index == 1853) return "H"  ;
    if (arc_index == 1897) return "W"  ;
    if (arc_index == 1905) return "W"  ;
    if (arc_index == 1923) return "E"  ;
    if (arc_index == 1936) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1940) return "H"  ;
    if (arc_index == 1946) return "E"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1949) return "E"  ;
    if (arc_index == 1952) return "E"  ;
    if (arc_index == 1953) return "E"  ;
    if (arc_index == 1954) return "E"  ;
    if (arc_index == 1969) return "W"  ;
    if (arc_index == 1987) return "W"  ;
    if (arc_index == 2001) return "W"  ;
    if (arc_index == 2013) return "E"  ;
    if (arc_index == 2023) return "E"  ;
    if (arc_index == 2024) return "E"  ;
    if (arc_index == 2034) return "E"  ;
    if (arc_index == 2035) return "E"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2040) return "E"  ;
    if (arc_index == 2043) return "E"  ;
    if (arc_index == 2066) return "H"  ;
    if (arc_index == 2122) return "W"  ;
    if (arc_index == 2170) return "W"  ;
    if (arc_index == 2171) return "W"  ;
    if (arc_index == 2177) return "H"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2224) return "E"  ;
    if (arc_index == 2247) return "H"  ;
    if (arc_index == 2300) return "H"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2421) return "E"  ;
    if (arc_index == 2422) return "H"  ;
    if (arc_index == 2434) return "H"  ;
    if (arc_index == 2442) return "H"  ;
    if (arc_index == 2460) return "H"  ;
    if (arc_index == 2469) return "W"  ;
    if (arc_index == 2475) return "W"  ;
    if (arc_index == 2477) return "E"  ;
    if (arc_index == 2483) return "E"  ;
    if (arc_index == 2485) return "E"  ;
    if (arc_index == 2486) return "E"  ;
    if (arc_index == 2508) return "E"  ;
    if (arc_index == 2516) return "E"  ;
    if (arc_index == 2540) return "E"  ;
    if (arc_index == 2557) return "E"  ;
    if (arc_index == 2566) return "E"  ;
    if (arc_index == 2589) return "E"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2619) return "H"  ;
    if (arc_index == 2662) return "H"  ;
    if (arc_index == 2670) return "E"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2685) return "E"  ;
    if (arc_index == 2686) return "E"  ;
    if (arc_index == 2687) return "E"  ;
    if (arc_index == 2688) return "W"  ;
    if (arc_index == 2689) return "E"  ;
    if (arc_index == 2690) return "E"  ;
    if (arc_index == 2691) return "E"  ;
    if (arc_index == 2692) return "E"  ;
    if (arc_index == 2693) return "E"  ;
    if (arc_index == 2694) return "E"  ;
    if (arc_index == 2695) return "W"  ;
    if (arc_index == 2696) return "E"  ;
    if (arc_index == 2697) return "E"  ;
    if (arc_index == 2698) return "E"  ;
    if (arc_index == 2699) return "W"  ;
    if (arc_index == 2700) return "E"  ;
    if (arc_index == 2701) return "W"  ;
    if (arc_index == 2702) return "W"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2704) return "E"  ;
    if (arc_index == 2705) return "E"  ;
    if (arc_index == 2713) return "E"  ;
    if (arc_index == 2717) return "H"  ;
    if (arc_index == 2755) return "H"  ;
    if (arc_index == 2762) return "H"  ;
    if (arc_index == 2770) return "H"  ;
    if (arc_index == 2793) return "H"  ;
    if (arc_index == 2803) return "H"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2842) return "E"  ;
    if (arc_index == 2854) return "E"  ;
    if (arc_index == 2856) return "E"  ;
    if (arc_index == 2860) return "E"  ;
    if (arc_index == 2861) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2881) return "E"  ;
    if (arc_index == 2903) return "W"  ;
  end 
  if ((thisRowAddr == 7) & (thisColAddr == 11)) begin 
    if (arc_index == 57) return "H"  ;
    if (arc_index == 146) return "H"  ;
    if (arc_index == 168) return "H"  ;
    if (arc_index == 234) return "H"  ;
    if (arc_index == 318) return "H"  ;
    if (arc_index == 427) return "H"  ;
    if (arc_index == 543) return "H"  ;
    if (arc_index == 566) return "H"  ;
    if (arc_index == 597) return "H"  ;
    if (arc_index == 632) return "H"  ;
    if (arc_index == 646) return "H"  ;
    if (arc_index == 711) return "H"  ;
    if (arc_index == 777) return "H"  ;
    if (arc_index == 930) return "H"  ;
    if (arc_index == 1034) return "H"  ;
    if (arc_index == 1038) return "H"  ;
    if (arc_index == 1048) return "H"  ;
    if (arc_index == 1049) return "H"  ;
    if (arc_index == 1050) return "H"  ;
    if (arc_index == 1051) return "W"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1054) return "W"  ;
    if (arc_index == 1488) return "W"  ;
    if (arc_index == 1540) return "W"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1561) return "W"  ;
    if (arc_index == 1573) return "W"  ;
    if (arc_index == 1579) return "H"  ;
    if (arc_index == 1681) return "H"  ;
    if (arc_index == 1734) return "H"  ;
    if (arc_index == 1809) return "H"  ;
    if (arc_index == 1867) return "H"  ;
    if (arc_index == 1875) return "H"  ;
    if (arc_index == 1962) return "H"  ;
    if (arc_index == 2073) return "H"  ;
    if (arc_index == 2078) return "H"  ;
    if (arc_index == 2088) return "H"  ;
    if (arc_index == 2199) return "H"  ;
    if (arc_index == 2269) return "H"  ;
    if (arc_index == 2378) return "H"  ;
    if (arc_index == 2388) return "H"  ;
    if (arc_index == 2396) return "H"  ;
    if (arc_index == 2444) return "H"  ;
    if (arc_index == 2618) return "H"  ;
    if (arc_index == 2621) return "W"  ;
    if (arc_index == 2641) return "H"  ;
    if (arc_index == 2642) return "H"  ;
    if (arc_index == 2643) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2651) return "W"  ;
    if (arc_index == 2653) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2658) return "W"  ;
    if (arc_index == 2684) return "H"  ;
    if (arc_index == 2706) return "W"  ;
    if (arc_index == 2707) return "W"  ;
    if (arc_index == 2708) return "W"  ;
    if (arc_index == 2709) return "W"  ;
    if (arc_index == 2710) return "W"  ;
    if (arc_index == 2711) return "W"  ;
    if (arc_index == 2712) return "W"  ;
    if (arc_index == 2713) return "W"  ;
    if (arc_index == 2714) return "W"  ;
    if (arc_index == 2715) return "W"  ;
    if (arc_index == 2716) return "W"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2718) return "W"  ;
    if (arc_index == 2719) return "W"  ;
    if (arc_index == 2720) return "W"  ;
    if (arc_index == 2721) return "W"  ;
    if (arc_index == 2722) return "W"  ;
    if (arc_index == 2723) return "W"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2725) return "W"  ;
    if (arc_index == 2726) return "W"  ;
    if (arc_index == 2727) return "W"  ;
    if (arc_index == 2739) return "H"  ;
    if (arc_index == 2784) return "H"  ;
    if (arc_index == 2833) return "H"  ;
    if (arc_index == 2917) return "H"  ;
    if (arc_index == 2921) return "W"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 1)) begin 
    if (arc_index == 12) return "W"  ;
    if (arc_index == 79) return "H"  ;
    if (arc_index == 211) return "W"  ;
    if (arc_index == 256) return "H"  ;
    if (arc_index == 340) return "H"  ;
    if (arc_index == 389) return "H"  ;
    if (arc_index == 449) return "H"  ;
    if (arc_index == 472) return "W"  ;
    if (arc_index == 478) return "W"  ;
    if (arc_index == 492) return "W"  ;
    if (arc_index == 493) return "E"  ;
    if (arc_index == 565) return "H"  ;
    if (arc_index == 654) return "H"  ;
    if (arc_index == 668) return "H"  ;
    if (arc_index == 697) return "W"  ;
    if (arc_index == 773) return "W"  ;
    if (arc_index == 799) return "H"  ;
    if (arc_index == 952) return "H"  ;
    if (arc_index == 1601) return "H"  ;
    if (arc_index == 1756) return "H"  ;
    if (arc_index == 1808) return "H"  ;
    if (arc_index == 1888) return "W"  ;
    if (arc_index == 1889) return "H"  ;
    if (arc_index == 1897) return "H"  ;
    if (arc_index == 1934) return "H"  ;
    if (arc_index == 1984) return "H"  ;
    if (arc_index == 2029) return "W"  ;
    if (arc_index == 2110) return "H"  ;
    if (arc_index == 2115) return "H"  ;
    if (arc_index == 2221) return "H"  ;
    if (arc_index == 2232) return "E"  ;
    if (arc_index == 2291) return "H"  ;
    if (arc_index == 2353) return "W"  ;
    if (arc_index == 2466) return "H"  ;
    if (arc_index == 2552) return "H"  ;
    if (arc_index == 2555) return "H"  ;
    if (arc_index == 2556) return "H"  ;
    if (arc_index == 2557) return "H"  ;
    if (arc_index == 2561) return "H"  ;
    if (arc_index == 2566) return "H"  ;
    if (arc_index == 2567) return "H"  ;
    if (arc_index == 2571) return "H"  ;
    if (arc_index == 2585) return "H"  ;
    if (arc_index == 2598) return "W"  ;
    if (arc_index == 2663) return "H"  ;
    if (arc_index == 2671) return "E"  ;
    if (arc_index == 2706) return "H"  ;
    if (arc_index == 2728) return "E"  ;
    if (arc_index == 2729) return "E"  ;
    if (arc_index == 2730) return "E"  ;
    if (arc_index == 2731) return "E"  ;
    if (arc_index == 2732) return "E"  ;
    if (arc_index == 2733) return "E"  ;
    if (arc_index == 2734) return "E"  ;
    if (arc_index == 2735) return "E"  ;
    if (arc_index == 2736) return "E"  ;
    if (arc_index == 2737) return "E"  ;
    if (arc_index == 2738) return "E"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2740) return "E"  ;
    if (arc_index == 2741) return "E"  ;
    if (arc_index == 2742) return "E"  ;
    if (arc_index == 2743) return "E"  ;
    if (arc_index == 2744) return "E"  ;
    if (arc_index == 2745) return "E"  ;
    if (arc_index == 2746) return "E"  ;
    if (arc_index == 2747) return "E"  ;
    if (arc_index == 2748) return "E"  ;
    if (arc_index == 2749) return "E"  ;
    if (arc_index == 2761) return "H"  ;
    if (arc_index == 2806) return "H"  ;
    if (arc_index == 2838) return "W"  ;
    if (arc_index == 2859) return "W"  ;
    if (arc_index == 2861) return "E"  ;
    if (arc_index == 2862) return "E"  ;
    if (arc_index == 2864) return "E"  ;
    if (arc_index == 2865) return "E"  ;
    if (arc_index == 2866) return "E"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2871) return "E"  ;
    if (arc_index == 2872) return "E"  ;
    if (arc_index == 2873) return "E"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2876) return "E"  ;
    if (arc_index == 2877) return "E"  ;
    if (arc_index == 2893) return "W"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 4)) begin 
    if (arc_index == 26) return "W"  ;
    if (arc_index == 51) return "W"  ;
    if (arc_index == 58) return "W"  ;
    if (arc_index == 86) return "W"  ;
    if (arc_index == 101) return "H"  ;
    if (arc_index == 123) return "H"  ;
    if (arc_index == 185) return "H"  ;
    if (arc_index == 202) return "W"  ;
    if (arc_index == 239) return "W"  ;
    if (arc_index == 241) return "W"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 278) return "H"  ;
    if (arc_index == 301) return "H"  ;
    if (arc_index == 310) return "H"  ;
    if (arc_index == 328) return "W"  ;
    if (arc_index == 362) return "H"  ;
    if (arc_index == 366) return "H"  ;
    if (arc_index == 442) return "E"  ;
    if (arc_index == 456) return "E"  ;
    if (arc_index == 470) return "E"  ;
    if (arc_index == 471) return "H"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 519) return "E"  ;
    if (arc_index == 535) return "E"  ;
    if (arc_index == 560) return "E"  ;
    if (arc_index == 571) return "W"  ;
    if (arc_index == 574) return "W"  ;
    if (arc_index == 577) return "E"  ;
    if (arc_index == 587) return "H"  ;
    if (arc_index == 609) return "H"  ;
    if (arc_index == 676) return "H"  ;
    if (arc_index == 690) return "H"  ;
    if (arc_index == 693) return "H"  ;
    if (arc_index == 719) return "H"  ;
    if (arc_index == 726) return "H"  ;
    if (arc_index == 744) return "W"  ;
    if (arc_index == 750) return "W"  ;
    if (arc_index == 752) return "W"  ;
    if (arc_index == 755) return "W"  ;
    if (arc_index == 759) return "W"  ;
    if (arc_index == 761) return "W"  ;
    if (arc_index == 767) return "W"  ;
    if (arc_index == 769) return "W"  ;
    if (arc_index == 775) return "W"  ;
    if (arc_index == 777) return "W"  ;
    if (arc_index == 810) return "E"  ;
    if (arc_index == 816) return "W"  ;
    if (arc_index == 821) return "H"  ;
    if (arc_index == 882) return "H"  ;
    if (arc_index == 883) return "E"  ;
    if (arc_index == 891) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 951) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 959) return "E"  ;
    if (arc_index == 967) return "E"  ;
    if (arc_index == 972) return "W"  ;
    if (arc_index == 974) return "H"  ;
    if (arc_index == 996) return "H"  ;
    if (arc_index == 1008) return "H"  ;
    if (arc_index == 1025) return "H"  ;
    if (arc_index == 1047) return "H"  ;
    if (arc_index == 1062) return "H"  ;
    if (arc_index == 1078) return "H"  ;
    if (arc_index == 1079) return "E"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1086) return "E"  ;
    if (arc_index == 1088) return "E"  ;
    if (arc_index == 1089) return "E"  ;
    if (arc_index == 1091) return "E"  ;
    if (arc_index == 1093) return "E"  ;
    if (arc_index == 1094) return "E"  ;
    if (arc_index == 1141) return "E"  ;
    if (arc_index == 1149) return "E"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1185) return "W"  ;
    if (arc_index == 1197) return "W"  ;
    if (arc_index == 1280) return "W"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1337) return "W"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1388) return "W"  ;
    if (arc_index == 1391) return "W"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1459) return "W"  ;
    if (arc_index == 1465) return "W"  ;
    if (arc_index == 1466) return "W"  ;
    if (arc_index == 1477) return "W"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1484) return "W"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1614) return "W"  ;
    if (arc_index == 1623) return "H"  ;
    if (arc_index == 1625) return "H"  ;
    if (arc_index == 1645) return "H"  ;
    if (arc_index == 1647) return "E"  ;
    if (arc_index == 1655) return "E"  ;
    if (arc_index == 1663) return "E"  ;
    if (arc_index == 1670) return "E"  ;
    if (arc_index == 1694) return "W"  ;
    if (arc_index == 1697) return "W"  ;
    if (arc_index == 1717) return "E"  ;
    if (arc_index == 1727) return "E"  ;
    if (arc_index == 1730) return "E"  ;
    if (arc_index == 1734) return "E"  ;
    if (arc_index == 1736) return "E"  ;
    if (arc_index == 1737) return "E"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1744) return "E"  ;
    if (arc_index == 1747) return "E"  ;
    if (arc_index == 1755) return "E"  ;
    if (arc_index == 1778) return "H"  ;
    if (arc_index == 1784) return "H"  ;
    if (arc_index == 1794) return "W"  ;
    if (arc_index == 1798) return "W"  ;
    if (arc_index == 1808) return "W"  ;
    if (arc_index == 1812) return "W"  ;
    if (arc_index == 1826) return "E"  ;
    if (arc_index == 1832) return "E"  ;
    if (arc_index == 1833) return "E"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1837) return "E"  ;
    if (arc_index == 1844) return "E"  ;
    if (arc_index == 1847) return "E"  ;
    if (arc_index == 1859) return "W"  ;
    if (arc_index == 1877) return "W"  ;
    if (arc_index == 1889) return "W"  ;
    if (arc_index == 1898) return "W"  ;
    if (arc_index == 1904) return "W"  ;
    if (arc_index == 1911) return "H"  ;
    if (arc_index == 1915) return "H"  ;
    if (arc_index == 1919) return "H"  ;
    if (arc_index == 1933) return "H"  ;
    if (arc_index == 1946) return "H"  ;
    if (arc_index == 1958) return "H"  ;
    if (arc_index == 1963) return "W"  ;
    if (arc_index == 1980) return "W"  ;
    if (arc_index == 1981) return "W"  ;
    if (arc_index == 1982) return "E"  ;
    if (arc_index == 1983) return "E"  ;
    if (arc_index == 1991) return "E"  ;
    if (arc_index == 1992) return "W"  ;
    if (arc_index == 1994) return "W"  ;
    if (arc_index == 1996) return "E"  ;
    if (arc_index == 1998) return "E"  ;
    if (arc_index == 2001) return "W"  ;
    if (arc_index == 2006) return "H"  ;
    if (arc_index == 2013) return "H"  ;
    if (arc_index == 2023) return "H"  ;
    if (arc_index == 2032) return "H"  ;
    if (arc_index == 2050) return "W"  ;
    if (arc_index == 2055) return "E"  ;
    if (arc_index == 2057) return "E"  ;
    if (arc_index == 2058) return "E"  ;
    if (arc_index == 2103) return "W"  ;
    if (arc_index == 2104) return "W"  ;
    if (arc_index == 2109) return "W"  ;
    if (arc_index == 2132) return "H"  ;
    if (arc_index == 2148) return "H"  ;
    if (arc_index == 2149) return "H"  ;
    if (arc_index == 2154) return "H"  ;
    if (arc_index == 2171) return "E"  ;
    if (arc_index == 2220) return "E"  ;
    if (arc_index == 2223) return "E"  ;
    if (arc_index == 2236) return "E"  ;
    if (arc_index == 2243) return "H"  ;
    if (arc_index == 2254) return "W"  ;
    if (arc_index == 2257) return "W"  ;
    if (arc_index == 2276) return "W"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2313) return "H"  ;
    if (arc_index == 2357) return "W"  ;
    if (arc_index == 2364) return "W"  ;
    if (arc_index == 2457) return "W"  ;
    if (arc_index == 2464) return "E"  ;
    if (arc_index == 2470) return "E"  ;
    if (arc_index == 2472) return "E"  ;
    if (arc_index == 2488) return "H"  ;
    if (arc_index == 2497) return "H"  ;
    if (arc_index == 2502) return "H"  ;
    if (arc_index == 2508) return "H"  ;
    if (arc_index == 2510) return "H"  ;
    if (arc_index == 2518) return "H"  ;
    if (arc_index == 2567) return "E"  ;
    if (arc_index == 2574) return "E"  ;
    if (arc_index == 2685) return "H"  ;
    if (arc_index == 2691) return "H"  ;
    if (arc_index == 2706) return "H"  ;
    if (arc_index == 2707) return "H"  ;
    if (arc_index == 2728) return "H"  ;
    if (arc_index == 2738) return "H"  ;
    if (arc_index == 2750) return "H"  ;
    if (arc_index == 2751) return "E"  ;
    if (arc_index == 2752) return "E"  ;
    if (arc_index == 2753) return "E"  ;
    if (arc_index == 2754) return "E"  ;
    if (arc_index == 2755) return "E"  ;
    if (arc_index == 2756) return "E"  ;
    if (arc_index == 2757) return "E"  ;
    if (arc_index == 2758) return "E"  ;
    if (arc_index == 2759) return "E"  ;
    if (arc_index == 2760) return "W"  ;
    if (arc_index == 2761) return "W"  ;
    if (arc_index == 2762) return "W"  ;
    if (arc_index == 2763) return "E"  ;
    if (arc_index == 2764) return "E"  ;
    if (arc_index == 2765) return "W"  ;
    if (arc_index == 2766) return "W"  ;
    if (arc_index == 2767) return "W"  ;
    if (arc_index == 2768) return "E"  ;
    if (arc_index == 2769) return "E"  ;
    if (arc_index == 2770) return "W"  ;
    if (arc_index == 2771) return "W"  ;
    if (arc_index == 2774) return "W"  ;
    if (arc_index == 2778) return "W"  ;
    if (arc_index == 2781) return "W"  ;
    if (arc_index == 2783) return "H"  ;
    if (arc_index == 2785) return "H"  ;
    if (arc_index == 2789) return "H"  ;
    if (arc_index == 2793) return "H"  ;
    if (arc_index == 2804) return "H"  ;
    if (arc_index == 2815) return "H"  ;
    if (arc_index == 2823) return "W"  ;
    if (arc_index == 2827) return "W"  ;
    if (arc_index == 2828) return "H"  ;
    if (arc_index == 2834) return "W"  ;
    if (arc_index == 2840) return "W"  ;
    if (arc_index == 2847) return "W"  ;
    if (arc_index == 2855) return "E"  ;
    if (arc_index == 2888) return "E"  ;
    if (arc_index == 2890) return "E"  ;
    if (arc_index == 2893) return "W"  ;
    if (arc_index == 2901) return "E"  ;
    if (arc_index == 2911) return "E"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 4)) begin 
    if (arc_index == 123) return "H"  ;
    if (arc_index == 164) return "W"  ;
    if (arc_index == 189) return "W"  ;
    if (arc_index == 263) return "W"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 300) return "H"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 384) return "H"  ;
    if (arc_index == 493) return "H"  ;
    if (arc_index == 559) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 565) return "W"  ;
    if (arc_index == 570) return "W"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 609) return "H"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 664) return "E"  ;
    if (arc_index == 698) return "H"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 712) return "H"  ;
    if (arc_index == 748) return "W"  ;
    if (arc_index == 764) return "W"  ;
    if (arc_index == 771) return "W"  ;
    if (arc_index == 772) return "W"  ;
    if (arc_index == 777) return "W"  ;
    if (arc_index == 780) return "W"  ;
    if (arc_index == 781) return "W"  ;
    if (arc_index == 782) return "W"  ;
    if (arc_index == 784) return "W"  ;
    if (arc_index == 788) return "E"  ;
    if (arc_index == 790) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 843) return "H"  ;
    if (arc_index == 950) return "E"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 996) return "H"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1062) return "W"  ;
    if (arc_index == 1197) return "E"  ;
    if (arc_index == 1417) return "W"  ;
    if (arc_index == 1418) return "W"  ;
    if (arc_index == 1424) return "W"  ;
    if (arc_index == 1425) return "W"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1629) return "E"  ;
    if (arc_index == 1645) return "H"  ;
    if (arc_index == 1706) return "W"  ;
    if (arc_index == 1709) return "W"  ;
    if (arc_index == 1711) return "W"  ;
    if (arc_index == 1712) return "W"  ;
    if (arc_index == 1713) return "W"  ;
    if (arc_index == 1715) return "W"  ;
    if (arc_index == 1727) return "E"  ;
    if (arc_index == 1762) return "E"  ;
    if (arc_index == 1767) return "W"  ;
    if (arc_index == 1771) return "W"  ;
    if (arc_index == 1800) return "H"  ;
    if (arc_index == 1866) return "W"  ;
    if (arc_index == 1933) return "H"  ;
    if (arc_index == 1941) return "H"  ;
    if (arc_index == 1946) return "E"  ;
    if (arc_index == 1999) return "W"  ;
    if (arc_index == 2028) return "H"  ;
    if (arc_index == 2037) return "E"  ;
    if (arc_index == 2094) return "W"  ;
    if (arc_index == 2102) return "W"  ;
    if (arc_index == 2110) return "W"  ;
    if (arc_index == 2148) return "E"  ;
    if (arc_index == 2154) return "H"  ;
    if (arc_index == 2220) return "W"  ;
    if (arc_index == 2232) return "E"  ;
    if (arc_index == 2265) return "H"  ;
    if (arc_index == 2290) return "W"  ;
    if (arc_index == 2331) return "W"  ;
    if (arc_index == 2335) return "H"  ;
    if (arc_index == 2401) return "W"  ;
    if (arc_index == 2457) return "E"  ;
    if (arc_index == 2487) return "W"  ;
    if (arc_index == 2510) return "H"  ;
    if (arc_index == 2530) return "W"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2554) return "E"  ;
    if (arc_index == 2558) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2560) return "E"  ;
    if (arc_index == 2563) return "E"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2691) return "E"  ;
    if (arc_index == 2707) return "H"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2737) return "E"  ;
    if (arc_index == 2750) return "H"  ;
    if (arc_index == 2772) return "W"  ;
    if (arc_index == 2773) return "W"  ;
    if (arc_index == 2774) return "W"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2776) return "E"  ;
    if (arc_index == 2777) return "E"  ;
    if (arc_index == 2778) return "E"  ;
    if (arc_index == 2779) return "E"  ;
    if (arc_index == 2780) return "E"  ;
    if (arc_index == 2781) return "E"  ;
    if (arc_index == 2782) return "E"  ;
    if (arc_index == 2783) return "E"  ;
    if (arc_index == 2784) return "E"  ;
    if (arc_index == 2785) return "E"  ;
    if (arc_index == 2786) return "E"  ;
    if (arc_index == 2787) return "E"  ;
    if (arc_index == 2788) return "E"  ;
    if (arc_index == 2789) return "E"  ;
    if (arc_index == 2790) return "E"  ;
    if (arc_index == 2791) return "E"  ;
    if (arc_index == 2792) return "W"  ;
    if (arc_index == 2793) return "W"  ;
    if (arc_index == 2805) return "H"  ;
    if (arc_index == 2816) return "W"  ;
    if (arc_index == 2829) return "W"  ;
    if (arc_index == 2839) return "W"  ;
    if (arc_index == 2843) return "W"  ;
    if (arc_index == 2844) return "E"  ;
    if (arc_index == 2845) return "E"  ;
    if (arc_index == 2846) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2849) return "E"  ;
    if (arc_index == 2850) return "H"  ;
    if (arc_index == 2852) return "H"  ;
    if (arc_index == 2853) return "E"  ;
    if (arc_index == 2855) return "E"  ;
    if (arc_index == 2858) return "E"  ;
    if (arc_index == 2916) return "W"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 1)) begin 
    if (arc_index == 79) return "W"  ;
    if (arc_index == 145) return "H"  ;
    if (arc_index == 322) return "H"  ;
    if (arc_index == 389) return "H"  ;
    if (arc_index == 406) return "H"  ;
    if (arc_index == 449) return "H"  ;
    if (arc_index == 450) return "E"  ;
    if (arc_index == 478) return "E"  ;
    if (arc_index == 486) return "E"  ;
    if (arc_index == 493) return "E"  ;
    if (arc_index == 508) return "E"  ;
    if (arc_index == 515) return "H"  ;
    if (arc_index == 585) return "E"  ;
    if (arc_index == 631) return "H"  ;
    if (arc_index == 654) return "H"  ;
    if (arc_index == 668) return "H"  ;
    if (arc_index == 720) return "H"  ;
    if (arc_index == 734) return "H"  ;
    if (arc_index == 773) return "H"  ;
    if (arc_index == 774) return "H"  ;
    if (arc_index == 783) return "H"  ;
    if (arc_index == 799) return "H"  ;
    if (arc_index == 849) return "W"  ;
    if (arc_index == 865) return "H"  ;
    if (arc_index == 881) return "W"  ;
    if (arc_index == 950) return "E"  ;
    if (arc_index == 952) return "E"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 1018) return "H"  ;
    if (arc_index == 1084) return "W"  ;
    if (arc_index == 1424) return "W"  ;
    if (arc_index == 1600) return "E"  ;
    if (arc_index == 1601) return "E"  ;
    if (arc_index == 1667) return "H"  ;
    if (arc_index == 1748) return "H"  ;
    if (arc_index == 1808) return "H"  ;
    if (arc_index == 1822) return "H"  ;
    if (arc_index == 1889) return "H"  ;
    if (arc_index == 1897) return "H"  ;
    if (arc_index == 1934) return "H"  ;
    if (arc_index == 1955) return "H"  ;
    if (arc_index == 1957) return "E"  ;
    if (arc_index == 1963) return "H"  ;
    if (arc_index == 2044) return "W"  ;
    if (arc_index == 2050) return "H"  ;
    if (arc_index == 2115) return "H"  ;
    if (arc_index == 2176) return "H"  ;
    if (arc_index == 2221) return "H"  ;
    if (arc_index == 2232) return "H"  ;
    if (arc_index == 2287) return "H"  ;
    if (arc_index == 2357) return "H"  ;
    if (arc_index == 2532) return "H"  ;
    if (arc_index == 2552) return "H"  ;
    if (arc_index == 2555) return "H"  ;
    if (arc_index == 2556) return "H"  ;
    if (arc_index == 2557) return "H"  ;
    if (arc_index == 2561) return "H"  ;
    if (arc_index == 2566) return "H"  ;
    if (arc_index == 2567) return "E"  ;
    if (arc_index == 2571) return "E"  ;
    if (arc_index == 2585) return "E"  ;
    if (arc_index == 2663) return "E"  ;
    if (arc_index == 2671) return "E"  ;
    if (arc_index == 2729) return "H"  ;
    if (arc_index == 2730) return "H"  ;
    if (arc_index == 2733) return "H"  ;
    if (arc_index == 2734) return "H"  ;
    if (arc_index == 2739) return "E"  ;
    if (arc_index == 2740) return "E"  ;
    if (arc_index == 2741) return "E"  ;
    if (arc_index == 2743) return "E"  ;
    if (arc_index == 2745) return "W"  ;
    if (arc_index == 2746) return "W"  ;
    if (arc_index == 2747) return "W"  ;
    if (arc_index == 2748) return "W"  ;
    if (arc_index == 2761) return "W"  ;
    if (arc_index == 2772) return "H"  ;
    if (arc_index == 2794) return "E"  ;
    if (arc_index == 2795) return "W"  ;
    if (arc_index == 2796) return "W"  ;
    if (arc_index == 2797) return "E"  ;
    if (arc_index == 2798) return "E"  ;
    if (arc_index == 2799) return "E"  ;
    if (arc_index == 2800) return "E"  ;
    if (arc_index == 2801) return "E"  ;
    if (arc_index == 2802) return "E"  ;
    if (arc_index == 2803) return "E"  ;
    if (arc_index == 2804) return "E"  ;
    if (arc_index == 2805) return "E"  ;
    if (arc_index == 2806) return "E"  ;
    if (arc_index == 2807) return "E"  ;
    if (arc_index == 2808) return "E"  ;
    if (arc_index == 2809) return "E"  ;
    if (arc_index == 2810) return "E"  ;
    if (arc_index == 2811) return "E"  ;
    if (arc_index == 2812) return "E"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2814) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2827) return "H"  ;
    if (arc_index == 2851) return "H"  ;
    if (arc_index == 2859) return "H"  ;
    if (arc_index == 2866) return "E"  ;
    if (arc_index == 2872) return "H"  ;
    if (arc_index == 2877) return "H"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 7)) begin 
    if (arc_index == 16) return "H"  ;
    if (arc_index == 30) return "E"  ;
    if (arc_index == 43) return "E"  ;
    if (arc_index == 70) return "E"  ;
    if (arc_index == 92) return "E"  ;
    if (arc_index == 95) return "E"  ;
    if (arc_index == 133) return "E"  ;
    if (arc_index == 167) return "H"  ;
    if (arc_index == 176) return "H"  ;
    if (arc_index == 189) return "H"  ;
    if (arc_index == 198) return "H"  ;
    if (arc_index == 201) return "H"  ;
    if (arc_index == 206) return "H"  ;
    if (arc_index == 209) return "H"  ;
    if (arc_index == 210) return "H"  ;
    if (arc_index == 217) return "H"  ;
    if (arc_index == 219) return "H"  ;
    if (arc_index == 257) return "H"  ;
    if (arc_index == 261) return "W"  ;
    if (arc_index == 276) return "W"  ;
    if (arc_index == 281) return "W"  ;
    if (arc_index == 288) return "W"  ;
    if (arc_index == 301) return "W"  ;
    if (arc_index == 310) return "W"  ;
    if (arc_index == 312) return "W"  ;
    if (arc_index == 315) return "W"  ;
    if (arc_index == 344) return "H"  ;
    if (arc_index == 359) return "H"  ;
    if (arc_index == 428) return "H"  ;
    if (arc_index == 433) return "E"  ;
    if (arc_index == 503) return "E"  ;
    if (arc_index == 511) return "E"  ;
    if (arc_index == 516) return "E"  ;
    if (arc_index == 537) return "H"  ;
    if (arc_index == 547) return "W"  ;
    if (arc_index == 554) return "W"  ;
    if (arc_index == 557) return "W"  ;
    if (arc_index == 561) return "W"  ;
    if (arc_index == 564) return "W"  ;
    if (arc_index == 601) return "W"  ;
    if (arc_index == 613) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 629) return "W"  ;
    if (arc_index == 634) return "W"  ;
    if (arc_index == 649) return "E"  ;
    if (arc_index == 652) return "E"  ;
    if (arc_index == 653) return "H"  ;
    if (arc_index == 686) return "H"  ;
    if (arc_index == 710) return "W"  ;
    if (arc_index == 719) return "W"  ;
    if (arc_index == 736) return "W"  ;
    if (arc_index == 742) return "H"  ;
    if (arc_index == 749) return "E"  ;
    if (arc_index == 756) return "H"  ;
    if (arc_index == 758) return "H"  ;
    if (arc_index == 815) return "W"  ;
    if (arc_index == 816) return "W"  ;
    if (arc_index == 819) return "W"  ;
    if (arc_index == 821) return "W"  ;
    if (arc_index == 822) return "W"  ;
    if (arc_index == 826) return "W"  ;
    if (arc_index == 831) return "W"  ;
    if (arc_index == 832) return "W"  ;
    if (arc_index == 841) return "W"  ;
    if (arc_index == 844) return "E"  ;
    if (arc_index == 856) return "E"  ;
    if (arc_index == 887) return "H"  ;
    if (arc_index == 892) return "E"  ;
    if (arc_index == 921) return "E"  ;
    if (arc_index == 955) return "E"  ;
    if (arc_index == 967) return "E"  ;
    if (arc_index == 981) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1040) return "H"  ;
    if (arc_index == 1050) return "H"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1064) return "W"  ;
    if (arc_index == 1070) return "E"  ;
    if (arc_index == 1076) return "W"  ;
    if (arc_index == 1080) return "E"  ;
    if (arc_index == 1088) return "E"  ;
    if (arc_index == 1091) return "E"  ;
    if (arc_index == 1108) return "E"  ;
    if (arc_index == 1141) return "W"  ;
    if (arc_index == 1157) return "W"  ;
    if (arc_index == 1161) return "W"  ;
    if (arc_index == 1195) return "W"  ;
    if (arc_index == 1236) return "W"  ;
    if (arc_index == 1257) return "W"  ;
    if (arc_index == 1313) return "W"  ;
    if (arc_index == 1316) return "W"  ;
    if (arc_index == 1321) return "W"  ;
    if (arc_index == 1345) return "W"  ;
    if (arc_index == 1348) return "W"  ;
    if (arc_index == 1349) return "W"  ;
    if (arc_index == 1350) return "W"  ;
    if (arc_index == 1355) return "W"  ;
    if (arc_index == 1358) return "W"  ;
    if (arc_index == 1359) return "W"  ;
    if (arc_index == 1362) return "W"  ;
    if (arc_index == 1374) return "W"  ;
    if (arc_index == 1379) return "W"  ;
    if (arc_index == 1399) return "W"  ;
    if (arc_index == 1404) return "E"  ;
    if (arc_index == 1410) return "E"  ;
    if (arc_index == 1421) return "E"  ;
    if (arc_index == 1427) return "E"  ;
    if (arc_index == 1449) return "E"  ;
    if (arc_index == 1452) return "E"  ;
    if (arc_index == 1460) return "E"  ;
    if (arc_index == 1461) return "E"  ;
    if (arc_index == 1476) return "E"  ;
    if (arc_index == 1477) return "W"  ;
    if (arc_index == 1478) return "W"  ;
    if (arc_index == 1481) return "W"  ;
    if (arc_index == 1483) return "W"  ;
    if (arc_index == 1484) return "W"  ;
    if (arc_index == 1485) return "W"  ;
    if (arc_index == 1486) return "W"  ;
    if (arc_index == 1492) return "W"  ;
    if (arc_index == 1494) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1544) return "W"  ;
    if (arc_index == 1653) return "E"  ;
    if (arc_index == 1666) return "E"  ;
    if (arc_index == 1689) return "H"  ;
    if (arc_index == 1739) return "H"  ;
    if (arc_index == 1751) return "E"  ;
    if (arc_index == 1764) return "E"  ;
    if (arc_index == 1778) return "W"  ;
    if (arc_index == 1791) return "E"  ;
    if (arc_index == 1796) return "E"  ;
    if (arc_index == 1797) return "E"  ;
    if (arc_index == 1811) return "E"  ;
    if (arc_index == 1816) return "E"  ;
    if (arc_index == 1832) return "E"  ;
    if (arc_index == 1836) return "E"  ;
    if (arc_index == 1837) return "E"  ;
    if (arc_index == 1844) return "H"  ;
    if (arc_index == 1851) return "H"  ;
    if (arc_index == 1852) return "E"  ;
    if (arc_index == 1928) return "E"  ;
    if (arc_index == 1932) return "E"  ;
    if (arc_index == 1958) return "W"  ;
    if (arc_index == 1959) return "W"  ;
    if (arc_index == 1963) return "W"  ;
    if (arc_index == 1971) return "W"  ;
    if (arc_index == 1977) return "H"  ;
    if (arc_index == 1978) return "E"  ;
    if (arc_index == 1985) return "H"  ;
    if (arc_index == 1989) return "E"  ;
    if (arc_index == 1991) return "E"  ;
    if (arc_index == 1995) return "E"  ;
    if (arc_index == 1996) return "E"  ;
    if (arc_index == 2000) return "E"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2072) return "H"  ;
    if (arc_index == 2090) return "H"  ;
    if (arc_index == 2091) return "W"  ;
    if (arc_index == 2095) return "W"  ;
    if (arc_index == 2103) return "W"  ;
    if (arc_index == 2123) return "W"  ;
    if (arc_index == 2159) return "E"  ;
    if (arc_index == 2168) return "E"  ;
    if (arc_index == 2198) return "H"  ;
    if (arc_index == 2215) return "H"  ;
    if (arc_index == 2266) return "H"  ;
    if (arc_index == 2285) return "H"  ;
    if (arc_index == 2287) return "W"  ;
    if (arc_index == 2288) return "W"  ;
    if (arc_index == 2292) return "W"  ;
    if (arc_index == 2294) return "W"  ;
    if (arc_index == 2296) return "W"  ;
    if (arc_index == 2299) return "W"  ;
    if (arc_index == 2303) return "W"  ;
    if (arc_index == 2306) return "W"  ;
    if (arc_index == 2307) return "W"  ;
    if (arc_index == 2308) return "W"  ;
    if (arc_index == 2309) return "H"  ;
    if (arc_index == 2321) return "H"  ;
    if (arc_index == 2342) return "H"  ;
    if (arc_index == 2346) return "W"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2350) return "W"  ;
    if (arc_index == 2364) return "W"  ;
    if (arc_index == 2366) return "W"  ;
    if (arc_index == 2379) return "H"  ;
    if (arc_index == 2401) return "H"  ;
    if (arc_index == 2424) return "E"  ;
    if (arc_index == 2470) return "E"  ;
    if (arc_index == 2476) return "E"  ;
    if (arc_index == 2482) return "E"  ;
    if (arc_index == 2484) return "E"  ;
    if (arc_index == 2490) return "E"  ;
    if (arc_index == 2492) return "E"  ;
    if (arc_index == 2496) return "E"  ;
    if (arc_index == 2503) return "E"  ;
    if (arc_index == 2538) return "E"  ;
    if (arc_index == 2554) return "H"  ;
    if (arc_index == 2567) return "H"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2605) return "E"  ;
    if (arc_index == 2611) return "W"  ;
    if (arc_index == 2634) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2751) return "H"  ;
    if (arc_index == 2753) return "E"  ;
    if (arc_index == 2768) return "E"  ;
    if (arc_index == 2769) return "E"  ;
    if (arc_index == 2775) return "E"  ;
    if (arc_index == 2776) return "E"  ;
    if (arc_index == 2794) return "H"  ;
    if (arc_index == 2810) return "H"  ;
    if (arc_index == 2816) return "H"  ;
    if (arc_index == 2817) return "H"  ;
    if (arc_index == 2818) return "E"  ;
    if (arc_index == 2819) return "E"  ;
    if (arc_index == 2820) return "E"  ;
    if (arc_index == 2821) return "E"  ;
    if (arc_index == 2822) return "E"  ;
    if (arc_index == 2823) return "W"  ;
    if (arc_index == 2824) return "W"  ;
    if (arc_index == 2825) return "W"  ;
    if (arc_index == 2826) return "W"  ;
    if (arc_index == 2827) return "W"  ;
    if (arc_index == 2828) return "W"  ;
    if (arc_index == 2829) return "W"  ;
    if (arc_index == 2830) return "E"  ;
    if (arc_index == 2831) return "E"  ;
    if (arc_index == 2832) return "E"  ;
    if (arc_index == 2833) return "E"  ;
    if (arc_index == 2834) return "W"  ;
    if (arc_index == 2835) return "W"  ;
    if (arc_index == 2836) return "E"  ;
    if (arc_index == 2837) return "E"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2849) return "H"  ;
    if (arc_index == 2855) return "H"  ;
    if (arc_index == 2882) return "E"  ;
    if (arc_index == 2894) return "H"  ;
    if (arc_index == 2901) return "E"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2918) return "W"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 3)) begin 
    if (arc_index == 26) return "W"  ;
    if (arc_index == 164) return "W"  ;
    if (arc_index == 189) return "H"  ;
    if (arc_index == 263) return "W"  ;
    if (arc_index == 273) return "W"  ;
    if (arc_index == 333) return "W"  ;
    if (arc_index == 366) return "H"  ;
    if (arc_index == 450) return "H"  ;
    if (arc_index == 559) return "H"  ;
    if (arc_index == 565) return "W"  ;
    if (arc_index == 583) return "E"  ;
    if (arc_index == 623) return "W"  ;
    if (arc_index == 675) return "H"  ;
    if (arc_index == 705) return "W"  ;
    if (arc_index == 748) return "W"  ;
    if (arc_index == 764) return "H"  ;
    if (arc_index == 771) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 775) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 778) return "H"  ;
    if (arc_index == 780) return "E"  ;
    if (arc_index == 781) return "E"  ;
    if (arc_index == 782) return "E"  ;
    if (arc_index == 784) return "E"  ;
    if (arc_index == 785) return "E"  ;
    if (arc_index == 788) return "E"  ;
    if (arc_index == 790) return "E"  ;
    if (arc_index == 791) return "E"  ;
    if (arc_index == 909) return "H"  ;
    if (arc_index == 963) return "E"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1062) return "H"  ;
    if (arc_index == 1308) return "W"  ;
    if (arc_index == 1417) return "W"  ;
    if (arc_index == 1418) return "W"  ;
    if (arc_index == 1425) return "W"  ;
    if (arc_index == 1580) return "W"  ;
    if (arc_index == 1706) return "W"  ;
    if (arc_index == 1711) return "H"  ;
    if (arc_index == 1712) return "H"  ;
    if (arc_index == 1713) return "W"  ;
    if (arc_index == 1767) return "W"  ;
    if (arc_index == 1866) return "H"  ;
    if (arc_index == 1941) return "E"  ;
    if (arc_index == 1999) return "H"  ;
    if (arc_index == 2007) return "H"  ;
    if (arc_index == 2028) return "E"  ;
    if (arc_index == 2037) return "E"  ;
    if (arc_index == 2045) return "W"  ;
    if (arc_index == 2094) return "H"  ;
    if (arc_index == 2110) return "W"  ;
    if (arc_index == 2220) return "H"  ;
    if (arc_index == 2232) return "E"  ;
    if (arc_index == 2290) return "W"  ;
    if (arc_index == 2331) return "H"  ;
    if (arc_index == 2401) return "H"  ;
    if (arc_index == 2487) return "W"  ;
    if (arc_index == 2530) return "W"  ;
    if (arc_index == 2553) return "E"  ;
    if (arc_index == 2554) return "E"  ;
    if (arc_index == 2558) return "E"  ;
    if (arc_index == 2559) return "E"  ;
    if (arc_index == 2560) return "E"  ;
    if (arc_index == 2563) return "E"  ;
    if (arc_index == 2565) return "E"  ;
    if (arc_index == 2570) return "E"  ;
    if (arc_index == 2572) return "E"  ;
    if (arc_index == 2573) return "E"  ;
    if (arc_index == 2576) return "H"  ;
    if (arc_index == 2630) return "W"  ;
    if (arc_index == 2724) return "W"  ;
    if (arc_index == 2737) return "E"  ;
    if (arc_index == 2772) return "E"  ;
    if (arc_index == 2773) return "H"  ;
    if (arc_index == 2792) return "H"  ;
    if (arc_index == 2816) return "H"  ;
    if (arc_index == 2829) return "W"  ;
    if (arc_index == 2838) return "W"  ;
    if (arc_index == 2839) return "E"  ;
    if (arc_index == 2840) return "E"  ;
    if (arc_index == 2841) return "E"  ;
    if (arc_index == 2842) return "E"  ;
    if (arc_index == 2843) return "E"  ;
    if (arc_index == 2844) return "E"  ;
    if (arc_index == 2845) return "E"  ;
    if (arc_index == 2846) return "E"  ;
    if (arc_index == 2847) return "E"  ;
    if (arc_index == 2848) return "E"  ;
    if (arc_index == 2849) return "E"  ;
    if (arc_index == 2850) return "E"  ;
    if (arc_index == 2851) return "W"  ;
    if (arc_index == 2852) return "E"  ;
    if (arc_index == 2853) return "E"  ;
    if (arc_index == 2854) return "E"  ;
    if (arc_index == 2855) return "E"  ;
    if (arc_index == 2856) return "E"  ;
    if (arc_index == 2857) return "W"  ;
    if (arc_index == 2858) return "E"  ;
    if (arc_index == 2859) return "W"  ;
    if (arc_index == 2871) return "H"  ;
    if (arc_index == 2916) return "H"  ;
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 0)) begin 
    if (arc_index == 12) return "H"  ;
    if (arc_index == 211) return "H"  ;
    if (arc_index == 388) return "H"  ;
    if (arc_index == 472) return "H"  ;
    if (arc_index == 492) return "E"  ;
    if (arc_index == 581) return "H"  ;
    if (arc_index == 697) return "H"  ;
    if (arc_index == 786) return "H"  ;
    if (arc_index == 800) return "H"  ;
    if (arc_index == 931) return "H"  ;
    if (arc_index == 1084) return "H"  ;
    if (arc_index == 1733) return "H"  ;
    if (arc_index == 1888) return "H"  ;
    if (arc_index == 2021) return "H"  ;
    if (arc_index == 2029) return "H"  ;
    if (arc_index == 2116) return "H"  ;
    if (arc_index == 2242) return "H"  ;
    if (arc_index == 2353) return "H"  ;
    if (arc_index == 2423) return "H"  ;
    if (arc_index == 2598) return "H"  ;
    if (arc_index == 2795) return "H"  ;
    if (arc_index == 2838) return "H"  ;
    if (arc_index == 2860) return "H"  ;
    if (arc_index == 2861) return "E"  ;
    if (arc_index == 2862) return "E"  ;
    if (arc_index == 2863) return "E"  ;
    if (arc_index == 2864) return "E"  ;
    if (arc_index == 2865) return "E"  ;
    if (arc_index == 2866) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2868) return "E"  ;
    if (arc_index == 2869) return "E"  ;
    if (arc_index == 2870) return "E"  ;
    if (arc_index == 2871) return "E"  ;
    if (arc_index == 2872) return "E"  ;
    if (arc_index == 2873) return "E"  ;
    if (arc_index == 2874) return "E"  ;
    if (arc_index == 2875) return "E"  ;
    if (arc_index == 2876) return "E"  ;
    if (arc_index == 2877) return "E"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2879) return "E"  ;
    if (arc_index == 2880) return "E"  ;
    if (arc_index == 2881) return "E"  ;
    if (arc_index == 2893) return "H"  ;
  end 
  if ((thisRowAddr == 5) & (thisColAddr == 4)) begin 
    if (arc_index == 7) return "W"  ;
    if (arc_index == 13) return "W"  ;
    if (arc_index == 18) return "W"  ;
    if (arc_index == 26) return "W"  ;
    if (arc_index == 28) return "W"  ;
    if (arc_index == 34) return "H"  ;
    if (arc_index == 51) return "H"  ;
    if (arc_index == 58) return "H"  ;
    if (arc_index == 70) return "H"  ;
    if (arc_index == 86) return "H"  ;
    if (arc_index == 101) return "H"  ;
    if (arc_index == 123) return "H"  ;
    if (arc_index == 136) return "H"  ;
    if (arc_index == 142) return "E"  ;
    if (arc_index == 158) return "W"  ;
    if (arc_index == 160) return "W"  ;
    if (arc_index == 162) return "W"  ;
    if (arc_index == 185) return "W"  ;
    if (arc_index == 212) return "W"  ;
    if (arc_index == 216) return "W"  ;
    if (arc_index == 233) return "H"  ;
    if (arc_index == 246) return "W"  ;
    if (arc_index == 296) return "W"  ;
    if (arc_index == 309) return "W"  ;
    if (arc_index == 334) return "W"  ;
    if (arc_index == 362) return "W"  ;
    if (arc_index == 366) return "W"  ;
    if (arc_index == 373) return "W"  ;
    if (arc_index == 410) return "H"  ;
    if (arc_index == 439) return "H"  ;
    if (arc_index == 442) return "H"  ;
    if (arc_index == 454) return "E"  ;
    if (arc_index == 456) return "E"  ;
    if (arc_index == 475) return "E"  ;
    if (arc_index == 482) return "E"  ;
    if (arc_index == 494) return "H"  ;
    if (arc_index == 506) return "H"  ;
    if (arc_index == 510) return "E"  ;
    if (arc_index == 535) return "E"  ;
    if (arc_index == 553) return "W"  ;
    if (arc_index == 560) return "W"  ;
    if (arc_index == 572) return "E"  ;
    if (arc_index == 590) return "E"  ;
    if (arc_index == 602) return "W"  ;
    if (arc_index == 603) return "H"  ;
    if (arc_index == 610) return "W"  ;
    if (arc_index == 612) return "W"  ;
    if (arc_index == 624) return "W"  ;
    if (arc_index == 654) return "W"  ;
    if (arc_index == 656) return "W"  ;
    if (arc_index == 676) return "W"  ;
    if (arc_index == 693) return "W"  ;
    if (arc_index == 717) return "W"  ;
    if (arc_index == 719) return "H"  ;
    if (arc_index == 726) return "H"  ;
    if (arc_index == 745) return "W"  ;
    if (arc_index == 752) return "W"  ;
    if (arc_index == 769) return "E"  ;
    if (arc_index == 777) return "E"  ;
    if (arc_index == 785) return "E"  ;
    if (arc_index == 808) return "H"  ;
    if (arc_index == 822) return "H"  ;
    if (arc_index == 862) return "H"  ;
    if (arc_index == 890) return "H"  ;
    if (arc_index == 891) return "H"  ;
    if (arc_index == 896) return "H"  ;
    if (arc_index == 898) return "E"  ;
    if (arc_index == 943) return "E"  ;
    if (arc_index == 945) return "E"  ;
    if (arc_index == 953) return "H"  ;
    if (arc_index == 954) return "E"  ;
    if (arc_index == 972) return "E"  ;
    if (arc_index == 974) return "E"  ;
    if (arc_index == 988) return "E"  ;
    if (arc_index == 996) return "E"  ;
    if (arc_index == 1004) return "E"  ;
    if (arc_index == 1005) return "E"  ;
    if (arc_index == 1008) return "E"  ;
    if (arc_index == 1009) return "E"  ;
    if (arc_index == 1016) return "E"  ;
    if (arc_index == 1025) return "E"  ;
    if (arc_index == 1044) return "W"  ;
    if (arc_index == 1047) return "W"  ;
    if (arc_index == 1063) return "W"  ;
    if (arc_index == 1068) return "W"  ;
    if (arc_index == 1075) return "W"  ;
    if (arc_index == 1077) return "W"  ;
    if (arc_index == 1085) return "E"  ;
    if (arc_index == 1106) return "H"  ;
    if (arc_index == 1121) return "W"  ;
    if (arc_index == 1147) return "W"  ;
    if (arc_index == 1169) return "W"  ;
    if (arc_index == 1170) return "W"  ;
    if (arc_index == 1185) return "W"  ;
    if (arc_index == 1190) return "W"  ;
    if (arc_index == 1197) return "W"  ;
    if (arc_index == 1220) return "E"  ;
    if (arc_index == 1230) return "E"  ;
    if (arc_index == 1279) return "W"  ;
    if (arc_index == 1280) return "W"  ;
    if (arc_index == 1296) return "W"  ;
    if (arc_index == 1319) return "W"  ;
    if (arc_index == 1322) return "W"  ;
    if (arc_index == 1356) return "W"  ;
    if (arc_index == 1390) return "W"  ;
    if (arc_index == 1412) return "W"  ;
    if (arc_index == 1423) return "W"  ;
    if (arc_index == 1428) return "W"  ;
    if (arc_index == 1429) return "W"  ;
    if (arc_index == 1459) return "W"  ;
    if (arc_index == 1495) return "W"  ;
    if (arc_index == 1511) return "W"  ;
    if (arc_index == 1517) return "W"  ;
    if (arc_index == 1557) return "W"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1591) return "E"  ;
    if (arc_index == 1594) return "E"  ;
    if (arc_index == 1595) return "E"  ;
    if (arc_index == 1597) return "E"  ;
    if (arc_index == 1606) return "W"  ;
    if (arc_index == 1607) return "E"  ;
    if (arc_index == 1608) return "E"  ;
    if (arc_index == 1609) return "E"  ;
    if (arc_index == 1611) return "E"  ;
    if (arc_index == 1615) return "E"  ;
    if (arc_index == 1617) return "W"  ;
    if (arc_index == 1621) return "E"  ;
    if (arc_index == 1626) return "E"  ;
    if (arc_index == 1627) return "E"  ;
    if (arc_index == 1630) return "E"  ;
    if (arc_index == 1632) return "E"  ;
    if (arc_index == 1635) return "E"  ;
    if (arc_index == 1638) return "E"  ;
    if (arc_index == 1641) return "E"  ;
    if (arc_index == 1645) return "E"  ;
    if (arc_index == 1646) return "E"  ;
    if (arc_index == 1648) return "E"  ;
    if (arc_index == 1668) return "E"  ;
    if (arc_index == 1674) return "W"  ;
    if (arc_index == 1684) return "W"  ;
    if (arc_index == 1697) return "W"  ;
    if (arc_index == 1731) return "W"  ;
    if (arc_index == 1741) return "E"  ;
    if (arc_index == 1750) return "E"  ;
    if (arc_index == 1755) return "H"  ;
    if (arc_index == 1759) return "E"  ;
    if (arc_index == 1776) return "E"  ;
    if (arc_index == 1784) return "E"  ;
    if (arc_index == 1795) return "W"  ;
    if (arc_index == 1823) return "W"  ;
    if (arc_index == 1827) return "E"  ;
    if (arc_index == 1857) return "E"  ;
    if (arc_index == 1883) return "E"  ;
    if (arc_index == 1894) return "E"  ;
    if (arc_index == 1897) return "W"  ;
    if (arc_index == 1899) return "W"  ;
    if (arc_index == 1905) return "W"  ;
    if (arc_index == 1910) return "H"  ;
    if (arc_index == 1916) return "E"  ;
    if (arc_index == 1922) return "E"  ;
    if (arc_index == 1923) return "E"  ;
    if (arc_index == 1936) return "E"  ;
    if (arc_index == 1939) return "E"  ;
    if (arc_index == 1946) return "E"  ;
    if (arc_index == 1948) return "E"  ;
    if (arc_index == 1952) return "E"  ;
    if (arc_index == 1953) return "E"  ;
    if (arc_index == 1954) return "E"  ;
    if (arc_index == 1969) return "W"  ;
    if (arc_index == 1980) return "W"  ;
    if (arc_index == 1981) return "W"  ;
    if (arc_index == 1983) return "W"  ;
    if (arc_index == 1998) return "W"  ;
    if (arc_index == 2006) return "W"  ;
    if (arc_index == 2012) return "E"  ;
    if (arc_index == 2013) return "E"  ;
    if (arc_index == 2032) return "E"  ;
    if (arc_index == 2036) return "E"  ;
    if (arc_index == 2039) return "E"  ;
    if (arc_index == 2042) return "E"  ;
    if (arc_index == 2043) return "H"  ;
    if (arc_index == 2049) return "E"  ;
    if (arc_index == 2050) return "E"  ;
    if (arc_index == 2051) return "H"  ;
    if (arc_index == 2053) return "E"  ;
    if (arc_index == 2055) return "E"  ;
    if (arc_index == 2057) return "E"  ;
    if (arc_index == 2058) return "E"  ;
    if (arc_index == 2059) return "E"  ;
    if (arc_index == 2060) return "E"  ;
    if (arc_index == 2065) return "E"  ;
    if (arc_index == 2109) return "E"  ;
    if (arc_index == 2122) return "W"  ;
    if (arc_index == 2138) return "H"  ;
    if (arc_index == 2144) return "H"  ;
    if (arc_index == 2148) return "H"  ;
    if (arc_index == 2149) return "H"  ;
    if (arc_index == 2152) return "H"  ;
    if (arc_index == 2154) return "H"  ;
    if (arc_index == 2160) return "E"  ;
    if (arc_index == 2191) return "W"  ;
    if (arc_index == 2224) return "W"  ;
    if (arc_index == 2236) return "W"  ;
    if (arc_index == 2243) return "W"  ;
    if (arc_index == 2247) return "W"  ;
    if (arc_index == 2253) return "W"  ;
    if (arc_index == 2264) return "H"  ;
    if (arc_index == 2276) return "H"  ;
    if (arc_index == 2300) return "W"  ;
    if (arc_index == 2347) return "W"  ;
    if (arc_index == 2375) return "H"  ;
    if (arc_index == 2384) return "H"  ;
    if (arc_index == 2390) return "W"  ;
    if (arc_index == 2391) return "W"  ;
    if (arc_index == 2399) return "W"  ;
    if (arc_index == 2421) return "E"  ;
    if (arc_index == 2424) return "E"  ;
    if (arc_index == 2429) return "E"  ;
    if (arc_index == 2445) return "H"  ;
    if (arc_index == 2457) return "H"  ;
    if (arc_index == 2458) return "H"  ;
    if (arc_index == 2477) return "H"  ;
    if (arc_index == 2486) return "W"  ;
    if (arc_index == 2508) return "W"  ;
    if (arc_index == 2510) return "W"  ;
    if (arc_index == 2518) return "W"  ;
    if (arc_index == 2519) return "W"  ;
    if (arc_index == 2535) return "W"  ;
    if (arc_index == 2541) return "W"  ;
    if (arc_index == 2574) return "W"  ;
    if (arc_index == 2607) return "W"  ;
    if (arc_index == 2620) return "H"  ;
    if (arc_index == 2659) return "H"  ;
    if (arc_index == 2664) return "E"  ;
    if (arc_index == 2670) return "E"  ;
    if (arc_index == 2684) return "E"  ;
    if (arc_index == 2685) return "E"  ;
    if (arc_index == 2686) return "E"  ;
    if (arc_index == 2687) return "E"  ;
    if (arc_index == 2689) return "E"  ;
    if (arc_index == 2690) return "E"  ;
    if (arc_index == 2691) return "E"  ;
    if (arc_index == 2693) return "E"  ;
    if (arc_index == 2696) return "E"  ;
    if (arc_index == 2698) return "E"  ;
    if (arc_index == 2700) return "E"  ;
    if (arc_index == 2703) return "E"  ;
    if (arc_index == 2705) return "E"  ;
    if (arc_index == 2706) return "E"  ;
    if (arc_index == 2717) return "W"  ;
    if (arc_index == 2752) return "W"  ;
    if (arc_index == 2755) return "W"  ;
    if (arc_index == 2774) return "W"  ;
    if (arc_index == 2781) return "W"  ;
    if (arc_index == 2785) return "W"  ;
    if (arc_index == 2789) return "W"  ;
    if (arc_index == 2804) return "W"  ;
    if (arc_index == 2809) return "W"  ;
    if (arc_index == 2813) return "E"  ;
    if (arc_index == 2815) return "E"  ;
    if (arc_index == 2817) return "H"  ;
    if (arc_index == 2860) return "H"  ;
    if (arc_index == 2861) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2882) return "E"  ;
    if (arc_index == 2883) return "E"  ;
    if (arc_index == 2884) return "E"  ;
    if (arc_index == 2885) return "E"  ;
    if (arc_index == 2886) return "E"  ;
    if (arc_index == 2887) return "E"  ;
    if (arc_index == 2888) return "E"  ;
    if (arc_index == 2889) return "E"  ;
    if (arc_index == 2890) return "E"  ;
    if (arc_index == 2891) return "E"  ;
    if (arc_index == 2892) return "E"  ;
    if (arc_index == 2893) return "E"  ;
    if (arc_index == 2894) return "E"  ;
    if (arc_index == 2895) return "E"  ;
    if (arc_index == 2896) return "E"  ;
    if (arc_index == 2897) return "E"  ;
    if (arc_index == 2898) return "E"  ;
    if (arc_index == 2899) return "E"  ;
    if (arc_index == 2900) return "E"  ;
    if (arc_index == 2901) return "E"  ;
    if (arc_index == 2902) return "E"  ;
    if (arc_index == 2903) return "W"  ;
    if (arc_index == 2915) return "H"  ;
  end 
  if ((thisRowAddr == 3) & (thisColAddr == 11)) begin 
    if (arc_index == 11) return "H"  ;
    if (arc_index == 56) return "H"  ;
    if (arc_index == 179) return "H"  ;
    if (arc_index == 255) return "H"  ;
    if (arc_index == 432) return "H"  ;
    if (arc_index == 516) return "H"  ;
    if (arc_index == 558) return "H"  ;
    if (arc_index == 594) return "H"  ;
    if (arc_index == 616) return "H"  ;
    if (arc_index == 620) return "H"  ;
    if (arc_index == 622) return "H"  ;
    if (arc_index == 625) return "H"  ;
    if (arc_index == 626) return "H"  ;
    if (arc_index == 630) return "H"  ;
    if (arc_index == 632) return "H"  ;
    if (arc_index == 636) return "H"  ;
    if (arc_index == 637) return "H"  ;
    if (arc_index == 709) return "H"  ;
    if (arc_index == 711) return "H"  ;
    if (arc_index == 741) return "H"  ;
    if (arc_index == 830) return "H"  ;
    if (arc_index == 844) return "H"  ;
    if (arc_index == 975) return "H"  ;
    if (arc_index == 1128) return "H"  ;
    if (arc_index == 1154) return "H"  ;
    if (arc_index == 1404) return "H"  ;
    if (arc_index == 1482) return "H"  ;
    if (arc_index == 1491) return "H"  ;
    if (arc_index == 1547) return "W"  ;
    if (arc_index == 1548) return "W"  ;
    if (arc_index == 1556) return "W"  ;
    if (arc_index == 1758) return "W"  ;
    if (arc_index == 1777) return "H"  ;
    if (arc_index == 1779) return "H"  ;
    if (arc_index == 1932) return "H"  ;
    if (arc_index == 2065) return "H"  ;
    if (arc_index == 2073) return "H"  ;
    if (arc_index == 2111) return "H"  ;
    if (arc_index == 2160) return "H"  ;
    if (arc_index == 2286) return "H"  ;
    if (arc_index == 2379) return "W"  ;
    if (arc_index == 2380) return "W"  ;
    if (arc_index == 2383) return "W"  ;
    if (arc_index == 2385) return "W"  ;
    if (arc_index == 2397) return "H"  ;
    if (arc_index == 2415) return "H"  ;
    if (arc_index == 2467) return "H"  ;
    if (arc_index == 2553) return "H"  ;
    if (arc_index == 2596) return "H"  ;
    if (arc_index == 2626) return "H"  ;
    if (arc_index == 2628) return "H"  ;
    if (arc_index == 2629) return "H"  ;
    if (arc_index == 2630) return "H"  ;
    if (arc_index == 2635) return "H"  ;
    if (arc_index == 2636) return "H"  ;
    if (arc_index == 2637) return "H"  ;
    if (arc_index == 2642) return "H"  ;
    if (arc_index == 2658) return "H"  ;
    if (arc_index == 2711) return "H"  ;
    if (arc_index == 2839) return "H"  ;
    if (arc_index == 2882) return "H"  ;
    if (arc_index == 2904) return "W"  ;
    if (arc_index == 2905) return "W"  ;
    if (arc_index == 2906) return "W"  ;
    if (arc_index == 2907) return "W"  ;
    if (arc_index == 2908) return "W"  ;
    if (arc_index == 2909) return "W"  ;
    if (arc_index == 2910) return "W"  ;
    if (arc_index == 2911) return "W"  ;
    if (arc_index == 2912) return "W"  ;
    if (arc_index == 2913) return "W"  ;
    if (arc_index == 2914) return "W"  ;
    if (arc_index == 2915) return "W"  ;
    if (arc_index == 2916) return "W"  ;
    if (arc_index == 2917) return "W"  ;
    if (arc_index == 2918) return "W"  ;
    if (arc_index == 2919) return "W"  ;
    if (arc_index == 2920) return "W"  ;
    if (arc_index == 2921) return "W"  ;
    if (arc_index == 2922) return "W"  ;
    if (arc_index == 2923) return "W"  ;
    if (arc_index == 2924) return "W"  ;
    if (arc_index == 2925) return "W"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 0)) begin 
    if (arc_index == 786) return "W"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 0)) begin 
  end 
  if ((thisRowAddr == 1) & (thisColAddr == 11)) begin 
    if (arc_index == 551) return "W"  ;
    if (arc_index == 621) return "W"  ;
    if (arc_index == 628) return "W"  ;
    if (arc_index == 633) return "W"  ;
    if (arc_index == 1777) return "W"  ;
    if (arc_index == 1779) return "W"  ;
    if (arc_index == 2910) return "W"  ;
  end 
  if ((thisRowAddr == 11) & (thisColAddr == 9)) begin 
    if (arc_index == 252) return "E"  ;
    if (arc_index == 289) return "W"  ;
    if (arc_index == 361) return "E"  ;
    if (arc_index == 435) return "E"  ;
    if (arc_index == 620) return "W"  ;
    if (arc_index == 680) return "W"  ;
    if (arc_index == 731) return "E"  ;
    if (arc_index == 861) return "E"  ;
    if (arc_index == 864) return "E"  ;
    if (arc_index == 871) return "E"  ;
    if (arc_index == 944) return "E"  ;
    if (arc_index == 1043) return "W"  ;
    if (arc_index == 1248) return "W"  ;
    if (arc_index == 1342) return "W"  ;
    if (arc_index == 1497) return "E"  ;
    if (arc_index == 1513) return "E"  ;
    if (arc_index == 1562) return "W"  ;
    if (arc_index == 1563) return "W"  ;
    if (arc_index == 1564) return "W"  ;
    if (arc_index == 1565) return "W"  ;
    if (arc_index == 1568) return "W"  ;
    if (arc_index == 1569) return "W"  ;
    if (arc_index == 1571) return "W"  ;
    if (arc_index == 1574) return "W"  ;
    if (arc_index == 1578) return "W"  ;
    if (arc_index == 1640) return "E"  ;
    if (arc_index == 1801) return "E"  ;
    if (arc_index == 1896) return "E"  ;
    if (arc_index == 2003) return "E"  ;
    if (arc_index == 2016) return "E"  ;
    if (arc_index == 2022) return "E"  ;
    if (arc_index == 2209) return "E"  ;
    if (arc_index == 2325) return "E"  ;
    if (arc_index == 2428) return "E"  ;
    if (arc_index == 2575) return "E"  ;
    if (arc_index == 2640) return "W"  ;
    if (arc_index == 2646) return "W"  ;
    if (arc_index == 2648) return "W"  ;
    if (arc_index == 2649) return "W"  ;
    if (arc_index == 2652) return "W"  ;
    if (arc_index == 2657) return "W"  ;
    if (arc_index == 2659) return "W"  ;
    if (arc_index == 2660) return "W"  ;
    if (arc_index == 2673) return "E"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 11)) begin 
    if (arc_index == 62) return "E"  ;
    if (arc_index == 168) return "E"  ;
    if (arc_index == 195) return "E"  ;
    if (arc_index == 203) return "E"  ;
    if (arc_index == 290) return "E"  ;
    if (arc_index == 427) return "E"  ;
    if (arc_index == 566) return "E"  ;
    if (arc_index == 580) return "E"  ;
    if (arc_index == 597) return "E"  ;
    if (arc_index == 711) return "E"  ;
    if (arc_index == 772) return "E"  ;
    if (arc_index == 969) return "E"  ;
    if (arc_index == 1034) return "E"  ;
    if (arc_index == 1037) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1042) return "W"  ;
    if (arc_index == 1048) return "W"  ;
    if (arc_index == 1049) return "W"  ;
    if (arc_index == 1050) return "W"  ;
    if (arc_index == 1051) return "W"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1053) return "W"  ;
    if (arc_index == 1054) return "W"  ;
    if (arc_index == 1067) return "W"  ;
    if (arc_index == 1112) return "W"  ;
    if (arc_index == 1488) return "W"  ;
    if (arc_index == 1540) return "W"  ;
    if (arc_index == 1573) return "W"  ;
    if (arc_index == 1579) return "W"  ;
    if (arc_index == 1681) return "W"  ;
    if (arc_index == 1797) return "W"  ;
    if (arc_index == 1809) return "W"  ;
    if (arc_index == 1886) return "W"  ;
    if (arc_index == 2133) return "W"  ;
    if (arc_index == 2378) return "W"  ;
    if (arc_index == 2396) return "W"  ;
    if (arc_index == 2618) return "W"  ;
    if (arc_index == 2641) return "W"  ;
    if (arc_index == 2642) return "W"  ;
    if (arc_index == 2643) return "W"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2651) return "W"  ;
    if (arc_index == 2653) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2658) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2718) return "W"  ;
    if (arc_index == 2726) return "W"  ;
    if (arc_index == 2833) return "W"  ;
    if (arc_index == 2917) return "W"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 10)) begin 
    if (arc_index == 314) return "W"  ;
    if (arc_index == 551) return "E"  ;
    if (arc_index == 628) return "W"  ;
    if (arc_index == 633) return "W"  ;
    if (arc_index == 1346) return "W"  ;
    if (arc_index == 1766) return "W"  ;
    if (arc_index == 1777) return "E"  ;
    if (arc_index == 1779) return "E"  ;
    if (arc_index == 2101) return "E"  ;
    if (arc_index == 2105) return "E"  ;
    if (arc_index == 2111) return "E"  ;
    if (arc_index == 2628) return "W"  ;
    if (arc_index == 2910) return "W"  ;
  end 
  if ((thisRowAddr == 10) & (thisColAddr == 0)) begin 
    if (arc_index == 500) return "E"  ;
  end 
  if ((thisRowAddr == 9) & (thisColAddr == 0)) begin 
    if (arc_index == 383) return "E"  ;
    if (arc_index == 500) return "E"  ;
    if (arc_index == 505) return "E"  ;
    if (arc_index == 586) return "E"  ;
    if (arc_index == 947) return "E"  ;
    if (arc_index == 1022) return "E"  ;
    if (arc_index == 1526) return "E"  ;
    if (arc_index == 1536) return "E"  ;
    if (arc_index == 2515) return "E"  ;
    if (arc_index == 2581) return "E"  ;
  end 
  if ((thisRowAddr == 2) & (thisColAddr == 0)) begin 
    if (arc_index == 388) return "E"  ;
    if (arc_index == 492) return "E"  ;
    if (arc_index == 581) return "E"  ;
    if (arc_index == 800) return "E"  ;
    if (arc_index == 849) return "E"  ;
    if (arc_index == 881) return "E"  ;
    if (arc_index == 931) return "E"  ;
    if (arc_index == 1084) return "E"  ;
    if (arc_index == 1424) return "E"  ;
    if (arc_index == 1733) return "E"  ;
    if (arc_index == 2021) return "E"  ;
    if (arc_index == 2044) return "E"  ;
    if (arc_index == 2116) return "E"  ;
    if (arc_index == 2242) return "E"  ;
    if (arc_index == 2423) return "E"  ;
    if (arc_index == 2663) return "E"  ;
    if (arc_index == 2671) return "E"  ;
    if (arc_index == 2745) return "E"  ;
    if (arc_index == 2795) return "E"  ;
    if (arc_index == 2860) return "E"  ;
    if (arc_index == 2863) return "E"  ;
    if (arc_index == 2867) return "E"  ;
    if (arc_index == 2868) return "E"  ;
    if (arc_index == 2869) return "E"  ;
    if (arc_index == 2874) return "E"  ;
    if (arc_index == 2878) return "E"  ;
    if (arc_index == 2879) return "E"  ;
    if (arc_index == 2880) return "E"  ;
    if (arc_index == 2881) return "E"  ;
  end 
  if ((thisRowAddr == 0) & (thisColAddr == 11)) begin 
    if (arc_index == 551) return "E"  ;
    if (arc_index == 633) return "W"  ;
    if (arc_index == 1777) return "W"  ;
    if (arc_index == 1779) return "W"  ;
    if (arc_index == 2910) return "W"  ;
  end 
  if ((thisRowAddr == 8) & (thisColAddr == 11)) begin 
    if (arc_index == 62) return "W"  ;
    if (arc_index == 146) return "W"  ;
    if (arc_index == 168) return "W"  ;
    if (arc_index == 195) return "W"  ;
    if (arc_index == 203) return "W"  ;
    if (arc_index == 290) return "W"  ;
    if (arc_index == 427) return "W"  ;
    if (arc_index == 566) return "W"  ;
    if (arc_index == 580) return "W"  ;
    if (arc_index == 597) return "W"  ;
    if (arc_index == 711) return "W"  ;
    if (arc_index == 772) return "W"  ;
    if (arc_index == 969) return "W"  ;
    if (arc_index == 1034) return "W"  ;
    if (arc_index == 1038) return "W"  ;
    if (arc_index == 1042) return "W"  ;
    if (arc_index == 1048) return "W"  ;
    if (arc_index == 1049) return "W"  ;
    if (arc_index == 1050) return "W"  ;
    if (arc_index == 1051) return "W"  ;
    if (arc_index == 1052) return "W"  ;
    if (arc_index == 1054) return "W"  ;
    if (arc_index == 1067) return "W"  ;
    if (arc_index == 1112) return "W"  ;
    if (arc_index == 1488) return "W"  ;
    if (arc_index == 1540) return "W"  ;
    if (arc_index == 1550) return "W"  ;
    if (arc_index == 1573) return "W"  ;
    if (arc_index == 1579) return "W"  ;
    if (arc_index == 1681) return "W"  ;
    if (arc_index == 1797) return "W"  ;
    if (arc_index == 1809) return "W"  ;
    if (arc_index == 1886) return "W"  ;
    if (arc_index == 2133) return "W"  ;
    if (arc_index == 2378) return "W"  ;
    if (arc_index == 2388) return "W"  ;
    if (arc_index == 2396) return "W"  ;
    if (arc_index == 2618) return "W"  ;
    if (arc_index == 2641) return "W"  ;
    if (arc_index == 2642) return "W"  ;
    if (arc_index == 2643) return "W"  ;
    if (arc_index == 2644) return "W"  ;
    if (arc_index == 2645) return "W"  ;
    if (arc_index == 2647) return "W"  ;
    if (arc_index == 2651) return "W"  ;
    if (arc_index == 2653) return "W"  ;
    if (arc_index == 2656) return "W"  ;
    if (arc_index == 2658) return "W"  ;
    if (arc_index == 2661) return "W"  ;
    if (arc_index == 2715) return "W"  ;
    if (arc_index == 2718) return "W"  ;
    if (arc_index == 2726) return "W"  ;
    if (arc_index == 2833) return "W"  ;
    if (arc_index == 2917) return "W"  ;
  end 
endfunction


// This is device placement generated from the qap solver used before hardcoded in mcmf.py file right now  
function MeshID lookupNoCAddr(ProcID currProcId); 
  case (currProcId)
    0: return 66; 
    1: return 100; 
    2: return 88; 
    3: return 86; 
    4: return 115; 
    5: return 113; 
    6: return 136; 
    7: return 56; 
    8: return 106; 
    9: return 31; 
    10: return 92; 
    11: return 20; 
    12: return 68; 
    13: return 82; 
    14: return 34; 
    15: return 90; 
    16: return 126; 
    17: return 109; 
    18: return 137; 
    19: return 127; 
    20: return 85; 
    21: return 75; 
    22: return 84; 
    23: return 49; 
    24: return 93; 
    25: return 7; 
    26: return 48; 
    27: return 70; 
    28: return 35; 
    29: return 114; 
    30: return 135; 
    31: return 32; 
    32: return 22; 
    33: return 140; 
    34: return 16; 
    35: return 2; 
    36: return 122; 
    37: return 45; 
    38: return 30; 
    39: return 138; 
    40: return 26; 
    41: return 74; 
    42: return 110; 
    43: return 36; 
    44: return 101; 
    45: return 123; 
    46: return 133; 
    47: return 131; 
    48: return 67; 
    49: return 37; 
    50: return 54; 
    51: return 130; 
    52: return 58; 
    53: return 102; 
    54: return 98; 
    55: return 97; 
    56: return 117; 
    57: return 116; 
    58: return 103; 
    59: return 129; 
    60: return 69; 
    61: return 46; 
    62: return 139; 
    63: return 17; 
    64: return 6; 
    65: return 89; 
    66: return 18; 
    67: return 44; 
    68: return 125; 
    69: return 96; 
    70: return 83; 
    71: return 142; 
    72: return 60; 
    73: return 52; 
    74: return 62; 
    75: return 51; 
    76: return 80; 
    77: return 5; 
    78: return 38; 
    79: return 14; 
    80: return 9; 
    81: return 42; 
    82: return 55; 
    83: return 39; 
    84: return 53; 
    85: return 104; 
    86: return 65; 
    87: return 50; 
    88: return 61; 
    89: return 79; 
    90: return 28; 
    91: return 134; 
    92: return 15; 
    93: return 76; 
    94: return 118; 
    95: return 8; 
    96: return 77; 
    97: return 112; 
    98: return 87; 
    99: return 94; 
    100: return 128; 
    101: return 73; 
    102: return 78; 
    103: return 91; 
    104: return 19; 
    105: return 105; 
    106: return 33; 
    107: return 57; 
    108: return 71; 
    109: return 81; 
    110: return 99; 
    111: return 124; 
    112: return 27; 
    113: return 41; 
    114: return 111; 
    115: return 29; 
    116: return 1; 
    117: return 121; 
    118: return 21; 
    119: return 59; 
    120: return 143; 
    121: return 72; 
    122: return 63; 
    123: return 95; 
    124: return 13; 
    125: return 40; 
    126: return 4; 
    127: return 25; 
    128: return 43; 
    129: return 3; 
    130: return 12; 
    131: return 64; 
    132: return 47; 
  endcase 
endfunction 
